-- de0clock.vhd

-- Generated using ACDS version 21.1 842

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity de0clock is
	port (
		ref_clk_clk        : in  std_logic := '0'; --      ref_clk.clk
		ref_reset_reset    : in  std_logic := '0'; --    ref_reset.reset
		reset_source_reset : out std_logic;        -- reset_source.reset
		sdram_clk_clk      : out std_logic;        --    sdram_clk.clk
		sys_clk_clk        : out std_logic         --      sys_clk.clk
	);
end entity de0clock;

architecture rtl of de0clock is
	component de0clock_sys_sdram_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component de0clock_sys_sdram_pll_0;

begin

	sys_sdram_pll_0 : component de0clock_sys_sdram_pll_0
		port map (
			ref_clk_clk        => ref_clk_clk,        --      ref_clk.clk
			ref_reset_reset    => ref_reset_reset,    --    ref_reset.reset
			sys_clk_clk        => sys_clk_clk,        --      sys_clk.clk
			sdram_clk_clk      => sdram_clk_clk,      --    sdram_clk.clk
			reset_source_reset => reset_source_reset  -- reset_source.reset
		);

end architecture rtl; -- of de0clock
