��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��5�������B���8���"���FE�Ҧ�@�Q\_������C]���5��1)2���� hڻ%pj�j��m���4 �w����4��O��� �P�˛����+���r\�8��s�;ۘ}�y���誛�I�e����-a�j��,C*��������~���>��75p�KcL�]�r��oՌ�I��r뎌 (��,H�grJ0�l���C-v��)���d�GFZ�bjU�zȱ%T��}X��?��~^u7�F�����ԝV�@:�2�9)�T�[���T+!w%�A����E��Eg�UWe���N�Aq�w2��>�;�b|c�������u#��W�R?�� �-��Fx��1�o�U���̈QU�_~�\�k���4��OAܥ(����GK>E�� 6�|M��:�GEO��d�[�	�_%��(%��S�S��[�ڔ������	r!qY>��'���7l�~ODǬ	s��MM�-!q�G,���d~w^j%�������w�j�|�ejF?k�3�R�x��J���?�BPU#�aT����	���8����~oD �Mz���y�w�]�o�U����[N�-�>aH0$��#�\��@SS�o5_�Q��[i��e��l~��8e��q-���/G;/*���P4��V���a��F<�T��
���P�V4��,�I*뢻U��q"`��Y��cG�8��Mh�D7��"�Tqhs�6{���gn
(]MxF���#LϠ� l�@ڼ��x����5I+0��RN��AF�YB��8�# �d+a�,���
���wœ�zE ˣ�('�%��&����/e �-��T+A�܆I���Bs[\D���=$K�{���=4آ�%M�{�-���J�9[����3�0\�GN���%�]��š`)��죿�N�P��t�f~/M��bf��	P׽C��$��=f���	�û	�#���/S�D��R �2'�Aߡ\d[�\�F�����6�p��+�	�PP����3Հ�����8��5	�8�f>����L�*�ɏ#?+o���d�v؄�;�~%K��^��nh" l��XEa�=|�8F~�5�<2�UF4[�(� bqXD�n��s���IȽ_uI[,�EANp��y����3��p
c��X��e*Ό�����O���e�c	yG���jH����	h{>_-&0ǉ�vNB�&w���-c+R�L#�KJ�@��y�<�'�ѡ�GE45���I/���0
>>Ite=kS���2�|]a1�{���E��\��Xe�^G�d)����t���3,^��&��nk�t�1�V8�wa;�e�����^K���d��8��Oꬂ<�DX������>�a���
�� 4<6:ĉ���%�O��vA��7i��`E3H��L��=�.���d{�Ы	']3K�k��n��F\�u�䠫'�1��[�l���И��J�w�]�����v$=0���gñKa�}Y�U(�������K���� �n�����>ۜ,���@R�E�קj\����a6� a$��2�bH��Me�&�ݳ�^��hb/�_~Ш>Ӄ���P:7GkZ!'�e�� �G�+Ψ#�e���<�ID�IF����ʳ�'�=P��io�hC����O�-v����6|!3�_L�,�艧��S�3�D�OW��S���\j&�J��.@2C�4[�"�^32�wse�\H�Ղy��q�v9��2�1x4��ݕ2�O�#od��wb�p�^�f��f�>B��I�)Ex���v2*9�y: ��)p+T��ݬ0m",��7'�Ur�{��DE������{��g�S@�a�K$�o�2��d��^��74ݦ�%����� �^�7�����$,�4���x��}7r���5}��'�r��2*����rg�,Ӓ���p	�ƺsP�:ȯ�N^�@�W��;�����U%� ���'�Z�œ@-d�|^���>���@`�R"��B_Q���#w�QY��)���ʑ-���lĴ4��Sё��t}�ԣ0~X��!��H���C�M\���Yo�.K�E_�h���N�ck��>��sV+�v����XY �*��%�h��_=�s9
؀Dˠ���}��qm�áW�*��^�.][���I�[{�}��[���y���qC�zV˃�p��*�P�rê)�*<i���K�J[	��[�\/���j�;Q�B�Ҿ�c�:<N��*�A��/�!x<(a� ��Wy�k������?�%+"�u'U�;S�BЮ�}q�5�]9�v��!�=����ΰ���c '4H�~^�a�C�u���5#�?��?��X�; �6��~�\��+���{�al\�d�X'���Vg�8�.Q,o�n_j+�k����:u��\ǿ��9�Q�2<' �܏q�P�ٮ�ժ�,��$������]b��"�OSg�a!Q��4a{�>>Ge"�*(-K���f�Xo�<|`L�4�iAҔ%�P����F/"^z���i�gF�P	*�QK���;����
�-��tຼ2����]�^P�E�ӡժxnP^���%�k�)�׻z�gqe�N<��\�?�����!*���ީ�r��5+I����j�YC�����)�	os'D����]Z�Kԙ��.�#E���FB����5�A��L������2_���.��V��G S�Lk4��`Ȫ�M����a&G�#5 U��C��Z7����G�A��v�O���W����c�����Z�~\[���	Et��Ee��O��/�''w��TϪ3V����5���5���^����`[4��{�WZ�R��ں*!@Bz�h�4��8ڝ��I�"�G2�T��w���ԡ�%���M��������2?���i�q.4s1AT��%������Vʠ>�;�5�hM'6`�I}q/��0�!*W����Lc���KG�@�����1zy��8jw�e�_�)������]�ZR�n?M~�}v�(�^�r��~]6y�
���iښ݂����0�]��%�w���,7��s���	o>L_n��ߝ��}��2
�>�O�h�gD(�\d�s�q�&��O�lpt�a�=L	���r��AEQ͒#_���f�+{+��߿zZ��}w���;]�y�	�i�p\g�Z������uL}+֔�eސ���x� ��sE3���m�N�R�X�P�F��gu{�*i緿Z��͜��ۘ�d�w�w0�sÓ�/��o&vC�&1=/�;q�Hob�𔒲Aԁ�8C;{�%�1-`iW}���mՖ��,�N���^�&�/�m��q(ל4�Tsn٫��]��k����az��@,�:�7�qWE�y͉y��)g�{��ʥ�+o����I^��ݖp.@�M��.�d���]�z:l�v�~���E�*t4��j�:���d������>�f7J�6���Qm��A�����<[4	vt�����n�D����W�5n��_k��͡g)��hy�s�Z�g7Cӱ���t�jp�0���͹��#>³���N��&����:Kie-�86,�{	�N�8U�E�p,�FP�E`�!-`1����\e�O�T����_�̯�ܞ��.D�	1��l�L��Y�<�co���AI!�gJ�(�Ӄ�K���?B���M����]9��������#�<}��4wa���D��Ӏ3?MB�W��U�+t�!��5Fʃj|TQ��]��/w:NPk�u�^d���\���Ԉ�ݰIY�G�;�O9�|�]�AT�Z�7�!��x�ӷY�PM$���ki��2bSV�'�w���r'�`������`��b�W��;��:�;�����Gr@��2���)3��7�n������EøA��2]9��� �Jf7�5��-�����W�͓���wBr��0��Fm���}rhD�'�o8��\"x����9�����,+xw��7��9��l3�2�e+d�ۭ�7eY!ز�6U*i��<��4�F �ʬ��|�r:>B�G����`�+I��1$8�j{��.E�W4���������/�3y�0���/lD���&��P�=*��o^�o��x�N�� A�9��f��[����)4�mM��*��G��|6�7��]`m�x #(���ܸ�5K��'9�vcQ)��Ѓ�4j�>��?4��e��V���t�[Z�P�E���D��d���5��x� ե=6�G�\e�K>�j�I��7C�a�sp����
N���h�� c�0�����[��9����n��^�}�q�z���G������a�����gAk&NieN��8��_g�P�����`�B��#���) �l�b�HTStY����{�����f,��y^T�!Zxh�'���i0ܫ �C���d�L����\����o[��I��J岕��_�
�s������_�=hW�e�� .1[$$���l�l7\�	�{��)��_
u�	v�@�;>�7���N�N�o�U>������Q�T��n{�����cB�zI�q�Aʄ�o?����ծ#��o�A��\ �,��vjv�[~��o�+3_I[��۞���P:2�~?C ���V9؍c.��Q�l��<��X�w.�!����,J�'���|oL?	 �L��r�7Y+�}�ѸW_��{h�e�ʱ��<q����E�5g�̗���!��ӷF.~�И�t���1�ɚ��/�!�y��{k��Xf�����bX�y��=CAVsh8����y1���P� �i��j�uX�����J�L�WZX1(6B_�l6��)�W%t`�sRD���������7V�d���hAD��0���w�U|��g�
��.�J��rQ'�dT(d�c���k7�"F���/iX������AM?��yG?�4b�����Yl�cc6Yi�����w0��8���o���s�V�nN��#�-�)I�z��ĭWG}`^�=K5`I\����GT����pQ)�毬���]{�����T��U��G��Ƕ�+ʅ=���Ub�q��ia���n-���j�է	!��&��_�sVV�G�ˈl�i�S��@+dۅ��XW�R�R����g�}�%�����%��?'�,���d�x��2�K���@�E^�p}s�#���M>���������9c'"�fP����|��9mj���yw�j�`�(Q������S�!��}��A����� _��Te5Ojf&8�So������dW�ቿ�K��<�=��Y�^��u��տ:�U�[a;�|���<%���f���(��ٍ�y3VC�_�u>E��W$ٝ����O�#����9���=�@H�TO��\x���ף�7�臜/KI�J�Y W),�G�i:������ �)s�2��'3������
���֚
����L烑X��;�	���0�}�Er�oz۹�ƀ/,�ҹ�H
�F���!s핖��m{ Vw�*�jpC���@��QO�����H�(�a�#�����+����,���0��� �m�b��'�O@L�%Z���~��ߠt:�j_������6�B>���B�&�r�������0����::�n���	د��J�-�(Z����b����f���ʹ��
�a�y��?!�O`�K:���V����p��+��J�p��:/17��;zЙ�Yh O�2C�J��[a�5�A��!����|��m
�y����(���HJ�}d&��_�{���;��-!�����7�>�/���~FhS�l>^"氞���槊��(k
��"R�Z�D}�N����9���9�I'�
��z�y��6H�+�+ߪ�$5����Ud�B�U�+� t[�L��M��v���y~�x�[޻C�3�`E_1d�&ڳ����8�<�L�i�J��@�Cq��s�_Lo��6�10�$�l�hm�e&3ym~�4�������?z��B%��9a�e�(^FG��W};��8�L0g�'�5���5��C!�a?\g5�0�Կ�
�RRP��G�p���>���E����
^hF(]L�SY{J59�d���/L����l}��|�`W�K�+0YW#:�L��ArN�'�!��[�f�oĿ�Yw�J1�_��w�6wm	�H�$ћѮ�)�
����#��0K�N^��O��{�Y50� qb� ��L���&��Ѱ��@K$2̈`F�
ߺ�Ȑ����Y7ym