��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D����gP�������������44��Pg��w�k�n�L�t�=�ʠ̲J�=�	�$tG�讧��p,��sC��Xu�_ S�	��mZK�qnu�*u"ǋ<�L*�2S���!��i�އh���
������)�=k��l��hx��I��} ���l��CaoK^G����F�HE���}�-���8���C��)�6v��q+���BɃ״��0�Ўl���Ax�`93Di�j�]��0x��uHo8ȁ�h�+���]�,L��uS��|�>5��9�8>�U̒ �|�o=���{�
'�[	��ԄgI.��Rs���Z�GݲB�_/h�_g�ˢGmYAa/E���,Ӥ`�΁b�d�@��+
��kz<ˤ(�w����0C݊��L87�C��������z��H�w��ڻJ�:>A��>I�B	�KW�-H��
 �ѶJ��;�\�16Ji�,�z}�:d�9E��_����Z���o-�[Ɯ��F$v�KG�%Z�:�oA4w�)[����:��z�X�o=B�e|�_2��ͰUSo����I#ظu��#x	oC}�v�%����KBU�2 p3 e�+�0ʝ��l�;$랉�A��t�h�?\�<��d"]���xuB�@3�{��e40/���GC��������ھΛ�HWR4��M�q��q��x�Gf�5�AW@{�-��LX�d��փ��Z�$�|�t��u�z(t�]7C�ua�Q�t��>l̘�9qaD���5:Ee��LsQ�����yEE������ ��B���+'�0����@x5^�(�uWD��j��
K��Q�0b�9x-�-=n.h�d�%��ʾ�~�H�;��zć(�}����?�v��f��f�T��ѵ�B�1�qR'1�G���"�XD[@;�:��}��D�Zsj�����s���A�$bg��DMYiP�Ϋ� `���
�6{c����ɔ�2�W���8��Vq��>C�?��6�7r��>o?2�>���
����q�{�w��	�N|���;n3�L4>����26�HQ
_z`�`�ck�L�~��z��K�è�N��=ß�yN�(+[Xz�tǾ���f�0��]˄�_0��L�|�o�Z+W��Ɔ�z�'�K��7ָ����:�Ӥ��還�]4�/J�M�=��n�iVG��J��>E���ӿ��S�T��G۸���}	�ɸi�݈֡9$�DQS�&�����Nw����ʤ�R�1���foh!ZhŊ޳�P�,]��LT�}��ɿ��#���m�{���Lw�^-y54q�/�߭��p��g�~�8���9_9l���)�>�1Y��[
k�����葰�ш�����U�s�)0���_V[���d�$/�_�5Ag�Н�!�Q_��/�ڕw��USB'��G�I�dG�&��hZ����mo�/��(��Y�@�@B}Rݤ�,���V@d��.�e��]���ر�����΋�.1^��|�n�]U� g0Dz&�#�8b� wQr(J(SKT5}�����
|�u��}s�ԥ�,�a
��[�8%z��K���jJ�=��\�c�tiSdr�ے ��:,����b���y���������cne[6|�p�'�\��d�Nki���P�n�T�ֹ����pv+q�[���Zbԏ�e�.zw�ߍ����F�����f����L���y���6���b�V���4�5���=�ҕ-G�~�E��-9dɯu7�Oe���� �AO�6����S�]��9=���0{[�|ӏ���ӲnۙC�Y:}�U1�+,�4o��fD����#�57�F�-}�����/־c�Fh���,��|��B>�
}�u���O���ug�B��m�C�	�k�X�����+��I)0��G|_Z�t|#kEsY��������g���I�撤řF����Ca�n�R��k��s���I�pG6yyA_���^��d"�mD���N��r�-|G������*��=Ts~��ߣ�8�c���)���RL�U0$��(\����5��n���xk�@���8ki:�W��C⨤�,U,_"���!*)G~dp����E.pv(ecZ�X|���%8`���ߒ��1�GD��Rq�$Z������S�p�r��`GH������)�nw,3��^7m�Z��Ax��4 ��w�c��M������u)D��>-�f�l���#��H��XE��e�=�w�:W%�p�p+HD�XD8W��O�zGUh窷���;��7տ��9Q��V��bft]�嗠�~�`��w�D��t7İ�8����p��f>�B�v׋1%7��f��8P���"���*v~�'k<�xh��nPŮ/�(S(D2=�����F3,�K����l�RC���:_|Qj��H��w5�3�G��?��:�>����[��a�,�<�l�+	�a�f�3�~p��6=zѦ(���iq�N�ȩ��p���{m	���yM.�A��Y6k<���]7�;���ôZE����"����aա��`� 	,;���؎�������j�kp�����������(����L&bˈ(�
Gl�����DI����h���[�GS)D�fmSD(7���Sx��*�/�'7�_��όuFfB�h�4��O��[h�H
B��r8����Fm������n5/}A���Ǟ�PqǢ���yQDW�fŴ�X��(�E&����4J��������%��aؖy���OQ�ROh��2�х��'{�O?���=��v_���j!�� �-�<�Lu��mZ��C��)D�P�Ȫq�HT��1�v�Z���O/kzZ�M��І�ˊ��Be�lff�{���3_�?gN�a��F�~,]=h#�.�^e ���O��8ޥ�-mw�>�~�K��*��C�RэN���B%��j��BB���g��	�&�,e���o�3�.#[H�;Y�k�%��yp�d��ͽ=M�<�S�yt}��$i�Ӭ�t���h��xP���q�+ɵ���C�����֋��Y0\X+V����WԬ�u�>C<���)z���5�[����a�� �7�~e�<_:řǎ��O�3��?ӽ�3m��x��5	7� BI��N�;����l���!d�G�p^FN�g�����M�Yo���١3�A�� �TRP�~�=��=��kh��P�w�۪�.wu",�GqW ��?bs������@f�J�	1�ޣ����c�!J��?��V�߂��7I`ЌŸ���Ԏ}#�=A���T�&��Q���(��M��ʩ����r���W+j^)��D��1�=k?i�n��02�� �b�s�P�/Ɋ�
�;[��ՙ����@���@��*W򨖂D�g�W�yg J��]�
,�8�.P���ZA�劏|��B���seJ~�{��Z��>�����Qy8Ac>ҎǳRˍp_|���0�F	���%��fǨ�I�_J�*5�4���J �.�L����z��˹Gh%��v�q ���ڰL�B�����su·�!�����J�.�~��UGv}:B���m��-�!��n�B�obJ?�l~��s4�� h���dv>�<h߅��{R۱�JS�FZ<��2��ط!��Q��%�RYT	Z(���̶u��Q1@�v�b�Su6��اV�%c 4.�+*���ff.3�|()Z���_+Od�J@��d�(�-.�A{�x��e5>��������?&R�Þ�L�]�Y�g�Q)�F�F�U�&N5O��[�n�#g)�î�[/�޼a��9Y	�\�Jz�l�s"��Z��4�Z������M��\.s�/V�'n��6�k|����k��.q�,��f:��( U�m�1�v�`>7���x�e�?��ID������g�|H���h�Ԗ�#7�U>C:Q��H�����8��yϬ��b0Y���>��/�V�?�e\���`sI���S�6��}�
�ZMrIU�Y�M\-�K��2O;��⭢l,jO`s0����3ޟKp� !4i���� �f�����Ei��o;q8���F��kR�W�O�Q�}������q'�N�r��o��^L������8ӡ26���q�"ڰ%m?�D����bf5�8Děn��.��p_����������g1��� �=;)�
p�;�Gp�TQF�&Բk����%�\t앰����>�*��}�շ���-CUp�]d9��u�L�],���Z �+�?0�W0�^�C[$��p,}��<2���Y7�n]8t�}X�*s��[�Τ��|�O��h�+��� w�w�1����W[��''�����W|;�i��N�Fa�$"���^�gA���r��ݬ���kAR����G)������q��9��1��H|t�ѭ��y�$#��'�=�1�4l������f/��M��ĵ׮�7 ���[z����E���\x;4b�r�֔���D�E�a*�j��/-�.�;�;�XQ�2x?LijR�5^V�n��Lf��mm�m�~5{������lp��5+@;�%�{`�|�q!��U*`ZX�KO��J�Y��2zau,ف���;/1u2ߺ �Z(��/m�	N�����1�F:n�6/BZ�PުU1s�uq��2z���q�s�=��{�3%hm��Xj�#���	�[y�Uϓv�$�p�����w��?k�J�I�'�ଡ�����6{�"�Ͻ��1$˟>_B2!8$ tp�e��ǒN�Ԋ�~�\c�3�[FT�Dj�4MW4�����+yBe�[��}KO�KR���t�G�W����}1tˎU���b�2
�a�n�6W59z��8�N����>1a�{�S���ЗBk�䰈�Bv,�E���(��n&�����=- �,H2J�AϤ�Az�j�8���D>�i�A"��֭���,�ۤ��0O�~�EC�J�Ʊ*����di��:�G�4�e�~!G�T^�|��R�'���U?�����m��ua�&-JX�_�`C�o�5��w����e$V��5͠P&�h�s�n���]H�|{��=(���:�k��64�|\����5��%��l�R�*e�hF���ǤX����6���ٞ홴�_�-��MN�Ẓv	��2�`u>�`�YǨ�ڜ�~�s���\�(]s�^i������tw�8���pd"ňR�<����7ݓ���6�*�!�4=�dg����������}h��dH�
��Mn����i�(�M)]�Q��z��YI�A�S;.�J�Yy%�؜�j&�����̆Q_��2��H��nX�ͽ��F�����������'��C\�hY��g�-h�����3:��ݮ��Y	��}jԢ��y��F�kNv��xߐ����i��]��"/ 뵳^C]���5I��С�Ct�:"^��y��i~j�T�#�bu/����Ѿ�L<��S�J;%��0󚶐�Ye���3-됥�Ctl�"�RB\H>��Z�:��p�����i���gh��o ���L^�:-Y+��u�!�`��23��1����T���rZ* e������&��s�w\�!�P���:��CQxc�
�/���,0�G-�E�`*��$9��xC���h|ۢx9)�JDC��%��&Cu��D��E'�P��Y�g]w��B��+%������	#1Q�h�\����f^r^/����@?5
ǂFf �aG�߱�.�T�|FVõ���gL����pm�6(�^���I�Q
;捨五��S�C��*A���ra����M��R|)��UV9�d�m;F�C�r��i�$H��0\��<��;�R3���әY�5Ptf�i�4����䐻�-��'�x���}ޯ���� X�h�H��X�|I�(��~M�50id�*�����h�&�j�`��8�^��tѓ� N'�6
܇��2r`�ކ���[�J�Ľ���[V�,�@2B�L8�O���3
���V����	�-�4"���ϓ�#+�܉���$�e��KIuP�A�`�->� ���$qA�b[?�bvn��w��zH���Y������B��eD��Ȍ/`��T�������̯}�W7- ��Ve���Od�ζ�g�%���ŭPASi���$�-o=�>��뇕��bp*�濋b�+�)���
է�h���Z��V����lީ�OC��t�1��ަ�Z�ޥv�)�o��������e�h�ayZ�i
t��� "�𽷒RF��n&�c,�i:�<�-�f���?��~3ZHx�Eb��-lDp�U ��A�yk+{e���{X׆K��>xH�#l5����Y(�T_��<V�{�A'l��?�c֪��xg�E��Ǻ�ux��[/����$%��,��Y6xOa��x��� x���I�����}\�����;$��1�|9�c��:N�O��3K^���\_�Mj�	���",���ܨ�8n�D���y�u��u�S��#�*P�2��� 6L���9#�;�M��RQ� tY�H$l��QcS�
���~$�'�*Z���倵o�$~�$<q��7���m%jEc�������L��� �s-k�UV!�Z�#ܛ����B�w�0bATyN7�Yi�}�KK�tl,]Xz��Ynhi�x�G�}�E�X���U~�(I��3�����ʙ�|>8.Me��K�c��,�r����"���,�u�!\�6�����
�XK��!X\N8',$-}í��,b�����Gtڻ�VeN������_zڭ;c��?,KsU	���/�N�)��x�7�ە9��0��U�Ɔ���xV��_�4�LY�<���
g$����O҄�M��8��k���G�,�S�����	P�o�EjW=��n@����sD��~ �z�g_��ϫ��(V�����Ž|�EY��_��(���)��ʉ����H;�a2���E9�|ֻ�!��p18ž��_r'P"D DiTӖ�DgԢ���s��K��q�O��FMa�7^륖� ��ն2Tq��\��27��t��s���w���bj�HA��t�+��S*+��3��_c$��2�SuE�@���*�rF�l�ō�y%ml߱
du���h�r�A��d�V�;���P��C�s[9r�hK ^�o��}@�L0���t���Z�,�dz�'C���F8����g��VRm�7��X��_���C��P.�4D[��0tM}\CZ�&�C�z���6�	�W���o��Ri\&慗@�=�A��!&� 	,p�b�zT��*�M]8k����a5È�˪����`��2,Y���閉�1n���q�����:���P�Ȥ�1����$V;j{qA���ݠ<��4];���7�@� �VM�)5D�0�ɽ[�
�����1�Iza�.8�'��0�|�p�'V�D�#���!%T�k�I���Gz���$c����ZϬ	-�FdC͐�7����36)�z�b����%�]y�n>p������������яh`w�>)6�^�S3�s���@ݗ��,*�;(�Xe���J��nQ�����>-+n��.��)�����Wy^s!��Ht�6� ݿ��ń�О��J�dm`:��Y���?21%TZb�d���"�7˞���1���x}l���D~����ڕ�ַ��-��W]�!�3��C���S��4(��[]���d�,474�O�xv���Y�S�~e
����{���N����"� ��&�m��&3�F��Q����G�Gp,�n���1�q����
}��qί��	k�FE�wS2�@��([윦2�>G���k�]�~`��Tآ�YɠKƑj+�s�j��U����g���>����|�_�MW���:D	z͙[��t.
j���Kʐ�#��0�6/�WH���z��'�S�zY�E��r�.�F��]����0�x!�98q�\��.4���T�o��ō���hC-�R���9$���BI
ū��`�h�;��B�,��D,fZ��>I|�e������;"�|Y�, ^)��	���#�2l��|��U�J��:�vTV�9Gmy�ĕ6y�s�3��</�&��W�D!��Ճ�bw�Tؑo[	5ҩ����޾��ٗcM��G��TP-�:n���?xs
l�-�_�eT��O]��˴P4 ����{+#x�S��+}�{a�Hf�	���Xh��R��O�ATI�?Az��R\le=������;�AŬ�_
P����K:�x�Ԓ��9'�1"�:���WR6�������@0E�r�AEjαu��̞�K[���|�1�C�,������d4��F!�/h�q��Hc3`\ T4,�2Av������cճ���}4ٟ1g3�I��67��3�;�]�v����yw84��w��<�y�* '���vۮ��o�e��iH�	"��6`|=Ĳ�9�M��> ziA��rn���Lޣ@�Y3Q�UO�d����+w��e#���9��;���E�s�����^�C��Q�#���Y�N�	�:� ��ye��(\���a&�G�6E嘵�g���5_m����\�SH�0v��B��dS�hס-bV�a�.��\C�s�lQ;q��:��)e�.�G�z�����zg^�~?98�o0�]�G�	�韀ǌ(�v���=J��
���?�~�����O�ErC&���G�[��5�άz���na���2s�V ���="L�{9�8�8��_�T|T�%��>�dҔ��{�`y�W�y	R�1�����N���%Gxi��&��{�»g�@��]!?t���L�պ@o(��Nݳ� p����=P���W3���܁2�#{��5��b+�t�>�p��T*h���O0�v-�	쳎�m7T�TM�p��zL0�6�d�a���Ҿ�����(�@�.����=�x_R	s�)��tu}k���*���E�BvJԃ���d:�g���+�U�wD�ߧu��bT��̄4�b��Ѿ��3h(��#��A�-�&yZh���1���Ê�.dдt�K����&���,[��;n<0�+��U�����_ѿ�]�r�=��뎈��t&�U�����i>%އs����b����}��9f�3 �q{�����Z���v� ��޾�Z���W��Ͽ�"�N�˳�o��W�մ�v0����n��~��ܶTz��.�E+�K3�UO1r�ݿ@%J��q��E�̈́��86ݑ���Xm����>��w�#k�ְ�P�_��3�$=K"��n�x�^�.�a@w�Y�����A��^� B�c�%_�Z��@e�6��b�V�܊^���W��<�8�Jl_E-�o�ڥ�AԦC}�;Voo*�m��3MA�j�(�Ғ"��A8 j9����͛�P(������\� �/�lv"�bg:X���FO�iˑk�������B���ɞu��"1��l7+.���e�|�yngU@�9m��rRl�!�w�7���Q�$.���U�ˆJ����F7�����xRi}-u�ƭ�U�����˵��X�ΜQ[J�'R����n��[04�a�bm����}��[9��w6p��`���o8b�#�d�n�v9��rdL�>�z1�FmY�z�H.�v�X��M�A׊B'�n�ǂ�e���3Y��;�u�[R��P,�\�?�wU����>_�@�W�s�_����o���_Pj����{��\Xe}�'?,6�q��n�E�|6�z�����O�\�h��1P���إ�o&�Lq��7e��O��y�l�* +�H}>���N�0��0_��h�c0$]�"qU�Ōn"h��߹)�{���k��!���Ι��,LN��� t�_���(+ͽ� ҽ�U�kR��"].��I��R������k8�H���\���=�����!"aZZ��_��ŊVR0�$
��A�)�L�I��",�;`'�h�����p97�/;W�O);a7<�౐K�����gFd�H�8�kB��}Yb��VI`.iŢ;���o��7NF���.=���sY�Y��E���k:]W�KzF�F 0���c�l�*/ݥ-'Br.���;ʜ�MerG�ĶohV)&��뭮�ٓ���}qY�ƚ�MڮJ�H8�:O}=�[u��
.�e�w�*9�
���_^�:(Ѿӻ�9v|�h�z5_C�}S2vw�����$�0L�T�)�	�á�7��,�ۯXn`���I &Zl���Wu��B����G� �`8���`G�9�m�4?O:$+5�y���	ù�w�֙gP2j�&���8��쫋�	��2
Qֿ��^�n[�4���dQI�{>���gN�&�zj�d{�P�o����Y��6�(?�n�!k�{EM��ZE!9��0"E,�?"p_|�`�L��"zд��Ԥ�>��d^�v4���O^�X�k�q��X'��=q3�C�G�uu��XbL�E��^D/�bYDL�ҿ���'�QB/�k5��}�Wt�&�`����A`�I&�!���爛B�3����� ��6�qB�������eջ�0%�%�m�@ ��Ĉ� ���2凓U&n�znL���#����k0�ћ i`n�^-�\E�Z'ޡ��L/޸�0�|3�!�-"��i9x�����g��D�-s��*���\�_��w8����j�ܵG��(�& �b�D޻�;�8gk�vR'Ȑ@�k��A�| �4yk�u{:�*�l�6�M��}���5�����#(�)kͼ���b�v�-�`K����2�2����nLB������������s瞕V;A~�&*M�Smxۉ��Y���K��5#���wr�Ed ���.X�ښ�M�E��k��7�@�n,�0i�%Z ��6����z?6����������o����<�d�����ȋR�y	�ɗ����e��-a���o�Y�O�/_�x�Uz��Q����-��`�De�SV����U<:�5���76���)�M,�k��5��l�٘��RT����Ov��&
�`f��������¡�٪�lx��s<��K�|"z���(ZΘ_jñ�6��e�j��	ч7mɭo�n[ĸ�̲E�cVz�t�����ژ^D�	�]�M'� 0�`B56)3{D���Q��9��0�ћƆ�Ğ��eV=7�䶜�)�-���%\��>*Tų
.��bK+3o�L� G'!�P<��U`�`���ߺ�Ur�)i� �8xZtT��F�H��1��BeyF#�y�?�D�k�%>���NA���d=6u�䆿S܈�t:��`:O�:,�EZ�E�+p�$ҥ�����Zd:� М����L����2a�O����@7����=�0#��j�T=�zS܀�'��_�i�ޝ�v#^�(pP(b9���-ɟ���u(�"�v���'n|�ۆ�RSښy�wQ�v1o"~f}K��l'�I��ÏZ�ōd�t��~f�U'��Z ߇�Z��)�>�����-��k�R]׎c�k�8//��G�.�Mq*-�����4����-]��3��c��X��/�C��~1�v}QĜ� .�߂�������ʹ��V XW�yԥ٤���8�Zۻ���q($�.e�|KK���%� �/��ȗį SY\�'*��R,(�Q�f�v�ɱ~��5�<	�K4���z�EB�Ē0#��ʵu�O�N`�[8���1�1d��^�����lD�y_u����b��WC�Ӟ��y�ۘ�2:��C 0�~g�l+�j�A9��S����f���<�B�v�7ٞ�^;�LZʊ!cvn~1o�y{��V�X�{�i�S~�L�c4��clA��g�!��ජ�Gد/y� ����%G��6 ����<mht�U���"5oʇ�Y��r��-TO_��ik�X���~�$�wEcZ2��杕��R��67}d{f5�}�
rH��T7w�^���ʊ�M��$+�g�5P-:���8��k4墼Z�=t�?�'{bq@�`捖�*���#�'��֛�o%
��w�B�^��*Ty�_1�B����Ӑ,�(�Gu�]��<��2��Tj�%^����WJ�ې�}ZckK-�Q����M��cL�b 5�O-��H]�@���{���n�����L	}ڞ�ч�-�v��~���	g f�(&VA��2}D����Z3��R�	|��ܒ�Vc�[g��!8� �y�	sc�Z�(��e����+A�qS��� Ԣ=��#�3��5�bV%��?��z���������a�+�rJ�8�r�*Ҹ6�h��i�NIۋ����y��o��C��I�3Nw�Ur�D(P��6c��_�wo�)B��雷�Y�%c��/�e���CV%���8���[.!�ɬ��	lnk���/�!���ԟT������u�p^�J�����6W�O��:}���uN f�����ƻ�z��F�q,�i�aYƟI�Ehc�,i�4F|;��A�����S��@�R`�u� U�rp?���<�{C��w��D/GȈ�	���z�eFխP���k��h	ژ�S�q��I��ʤ�x9�}��X�m$�:�f����m`��$@0�kj�P��%(;Zj�Ǣ`����lƼ��nNQq������h3����=��7�UV�ƛt����hT ��K���8�$m !F�����\���qkr���k
���*�*�9��k���7}�.�!�g^ �U�zf��Ո�����z��~�<�v��8�˳�s�)�V�fC��Y^�v��1�r(�_Xʭ�׭�wUE��c�zx]�y[��X�Vư��U�9ύ����v�hN����Pם7�K9�u����З����t>i��C�'Z��D�Ll�2o\YN�ZɄl��O+bX�|H0&f�M�F�Rc<1q�w�\����nR�br�,�4{ 1��7ug����A�I�&� ��;m��L���k�h
�U�mV�а-��z��M���]�r�36�=��	L�V���xE�n���f�j?}��A��K���[�_E��V�-�/D��5�?*�������Y$�ߺIoz��3��?:��،2q<�����n�\��l��!����SH�7��8,��&��$��Q�`���2|Vf�z��I�)h8)C�T��ǒf�jeG�<)�z����ش?H��&r&W��Kg,��a�#��ƹB�	��ɫ��$���
���`s�%�)^|�h
R���)�����[��I3mP�HN��"�I�[x����t�|�#�D?�*�	$��ϋ�kVy-���	�1���^�@�@ ,D&w�|n\(
&+UL�Ӛ?�\������� CIP����A|� �ɼ)<�N=(C��c��0���@��bKAs��\G���-��R�CRŭ��!�|���?Ϟ�K�a	�Vy�r40P|�5�a�Xz�w9m�~ރCu�"�N���Yo�pH�J(A�)}jV�쟷�� wt��xu�L�c! �=�&%���^�"R�h&8�m����c#�s�F�&\�C� mQk��p�.H�w�ύʚ�s�U�J ��l���r��G�0#���3-	5~>E��ȉTH���qWog�ER�:�������f�P
�ǁ�����஥�|�,9\���~���P�sh��k��^�d�͓^���s|-`�N-����s^ߕ]Z��+$
؏O~z,Ԇ�r��.�}��������m�!t��}�<]O�g����7z�M��lIy�g�|`��j�j��R�e�X��;T�5�V���~==>ce��"H:�n:�3]���|�T�=��)����n���^ue��ʽ��v�����ꬳ�:�&m����5G�_Y�WA��\�M)]�~�9/�ٶ(ҳ�g'׳y���)�,�=��_�)!���x���?s6@1��9���R�<�w3��o�l�ZgMx� ��&©���Ϸ������kZ=��l��^���ڪi5�/b�1�Mе���TVH�`,nĪ�d<sZ�HE�8�G�Va�"]�r��g�J��P�أ���'�Lw"bv��p"}|��\9�Z���U:�A��4P�G�4>�Q�n�@�.3�׍�%��B��Զ9���_�S�崎�4�}�F�h��i�cnL�@�]9@����/�Rxű?=�m�(�Ջ�S��2*��Z]Z0������҇�+V�7�8�h/�N�:��#.���e���%�v�9ׯ�'�J�w!��P>�j"��|�)R���=�g�l�+i�ZgOޒ�)��`�1,����~���Z*4���l�O�������{�Hf6�2��׊PC��/�U��7>������G���~��.D�m�������i�'�2��b�{xE|&8�G�D�}R���,��+�`�
˥���D�mڜ䐺���x0;<C0m!K�&j��jP[*���qW�(�m����#�1]�ڗ�v��X�8۽��(��<�Ԣ��~DԻ��kձ���M�:�~hZ}��a�CG�y�'���^�ͻ�~�b�ʂ��+P�Z��J������M��R�r����sV�F/f� �<�=��|��	�ĸA���<�cfH������XW
�}���mD��T+z8�X�6:b��-�?9 }VOEv?� k�z7v9;"k�� �G��a��Jl�/ ��r�L�d}	:&��	?Ʊ�N��<��l�f�G�,B,��m98�c���QB.�Kr�`.��s�>TRR�>L�J
�T�#C;nY�(�i�oVF��Ԙ籓���;�Y�p���ph������\�(E>\V��H���Rx6.�3{xS�6��C"����hKc�|���#h=��ս���0�}��CP!��)��� K|Ubwԉ(U��7�==��b��}��p�lpZv�ke�$��U"5� HH�5��\7������Q%�����L���N��U�^K��5���v���<����m�L��f���E{���sd�~8P�X��%����D��\���lY���w�0��fq#f3��,�t�����"��\)O��ٵH��/P��?���{Gh�.�r^"-X�����p�j��\�KK�}��@5x7^��W�L�2�IV����0C�nV�u�4x\[�3�ĭ�����v6U�X��}簐#A�ká>]��6-Au)��v]cj�Y���ڶn�nj:?) P�7I�O^xF��� ���Ƒ��{5�<Nh,�A�98 �y�T��F���i7�!s�I�z?�t-eUrϢ��~�	Yg�b���x�B�/�2oyv�ԀK�B�!܃����@*-rv�ʋG���a&#�4�\'$��� ޣe��}��#��tZT/AG���2o.�p�(a{�3�E��H���zkb�~.\h��u/Q��6I7�O�v�x��w*{��]���3؉�e�����F%�2���r���0��{�X����a=?��������61$�ne8%q�\3��$
�Ws�~����<��eE�������#����q�|����g����=�Aѡ���p ��g�&|Uq�;�h��%D�!jEhh/�q��-�(]pH9_�������� �@����QU�03�'Ƥ���H�$'5��w��v�xHq��?�_"E l�T.����7��8�םV��ʼ����s��F~e��m2��8��/��5�m��f0	�1��AL�0�7��uQ�����e��6�ڔ_�Cm������D7sX7 9IX4�ޣ���\�B�=�$�LS�
�Q��=�PkǨ"Ob�b�x����+��S��C�o+"��{�ĉ>A��]N�~�Q��
D�"&KZCj�E�B���m�@ K�����n�%"N�G��{�Hx0:Jl
6��
��/-��"	��t�m�U��N�ɌF�eK����te/�E��𢎨G��3,
MG�Bf��;ꅕf�$P;s�͗uU�l��Ux�f �8R��n1\%��~N/� Ѯ����O���h�3V/����#ǝw�m��!�d�9ukG�o�_�B�M�$�	8#�6	������9C"c�(���4s����(��g[R�O�&�OC��͈K�"kx�6Yq����';u?g�f�9�Di�:�x�K���P0�"�h۟�(O��5/��Nm��T?�Q@/�a�SE�!�P�hFu�#�v����'1�3=�	�sP,8�Gq@d�g΍8����H�5K�Y����F���T
�]��y8�<I�W͌�a����A��׸�X��-!�B�RDZJ@��L���ٔ��HRQh[+� ��#!�m`QcT�`�����9# �3]?��ն	3��E\��o�-}R��+"��<��}ܴ7�N���H�w�v��BL;��BDvyhĀ�դwc��rT���5�'�7l�	���۾�^�&����h�L�:c�����$�4-��c��a񽓴���ȷ���>Aw����1�=���`2��{%���`�p2� �>E%&]�5�FC1�i�g�rD-�1�a��rv[����[]�~���G�����0<�5�ڻ\@_���.i�P �@n�.#�Y�0��乫~���_��avS@�
�#B��o�N����L��%�F5�ƙ>
C'j���0���?�n��:x(�h�����dO����4��Wj;U/�^�Oj�޳D�s��ȗ⢡>|h�?+�z�����^;��q�	�fA�gg*�Ɨ�׃�s��ѻ��x�
L溿޻�yQ 9>5H� t_FƁA�o#QX����%5U� �G�Tc/ku�=�F<��wY��V�������6V2�+{���!�?��+��i'<����|��Lo�,�^?{x��,���&Y�}f,8���1Q�)�tZ�6��`K�Ct�5o�|�+ӫr�2��1Y���� �"��,������d	֏�4}rxs���l�#
'}�X��:&�0���իG�0��&`�ORq�d+�:�r���ls�p+s �G�>���(k|�'�q��B~�V� �� ��Rr��L!r{�g��N+VF��Ҕ��_*X��?.�0���������� ͵�߶�~U���)W���ͅ�ގ�j�y�I�Wp��Ze����' �r#�����$�h4������TkK���`"�I�v��g%%�l�"z'��	�����^	lr`Dv�M���|��.��f�x��"_7��5v������W�7s�����x�]���� E�D��+��Dx��ٵvG#�h�n�=��&|?C#�Y���~�ӻ�Ʒ&rȲ^ѤB�!�����Jx��{ �jh'"�D�oZ�������o�����AHez�u��U~
�/Z�a(�ɸ?x�v���'Σ��gL���$����J$�̏dG�o�$�ބ�!������A؋;���/5���ߦ�C#��Q�Cw.�"`Y��JFVR��Q�B��Ğ�����Ds�>��Z��||g�����XMy8�$�������7���\��<z+�V��ӽp��6�4W���2�[��;}��.ǓE�����p�����@�+XHY�q��e{�Y�h7H_4��O�1V@[^�OԪ󪁜�Ej�6K ����B�+w��:-�.��>q��	�D�42g�խ1*���;̡	�V8cIa4f���!�:kd�0SI\^m�v�?,K�Q�a����P"�3]R�=Z���+(G�t6�����t�/�{�P¦J���Ni�W^+�7�w�m���SϦ������7���'��Y�sG�����M9F���&k]�4S��~�ا�ˣk|����b�Ny��j&���=�tM��أѾ�o�p1~~r�o-��
}A('�m��]�$)iE�'�/�B�8����V��~��j��b:q���-�+WO��0�ZߜI?YCQt:v��/����#*2� i�}WF��i��_B��í��`���S#�Y /���3��0�>$���ԛ����j��A!�� �02�|�l(�.=����\G���,�F�\�iӌ�W���'���D�rn���(V��U4���q�Q<N5`�	�}ű�h#���{H,�F5ﳨ���Z�-�qF�w�����˂��J*侇Nr1��S ld�2xMc��" ���Hf��.x�����"���w0��^`H�bC��Os��c�)���Ȓig�k�p�\(I_]�]Q��y,sS*�N%,]86���.���vY�J���s����1T�<���݇L��-��5B�qD�;������]We��.%��!pgz<�G�'������?��>��G�#O�x�g1W�� �
�����း*��,�7�P�e�8f.��(tE�C3w��!������:r���{�f�F�,k�sތ���ciaʂ~����SRH��&β��^�e��D��
���v׷�&��Gn��o3���J���|��x���0N����bEn�4�dޒ���+L�!�����8� /�p��#�ǿP��BO��U����"ƘHT*�D�C�*BO��j��<���-r#=^}q(l&�m��3<� ڌ	VME�����Fu-�X���L#%l�������(s��r�[�j�2�8Phy�����t�@p3&��P~>�6�Om��6�꒏��9�+��}  /WqZ��2��dJG�[�A0�
d
�|�h�W����Jcz�p�;�m^��ıJ���((A�����D�f�9�� Er|<��ODA�O�R\�8p������?{�ۦS.ᚖ�O�r,S+B����	>Z"�sQ�i�[��Pȱ�p���X	%���Wڵx�1�������G�������Q��I+�Ι��oŉ��aa8<��d��F_����2�D��$��rE��b�O�z��d�S���*9�y�n:�y��`��¹������w�O�97��r�T���x�'}���w�
5�����y�&fr�胺�
+D�N�
v}�o�ؠ�x���Y��ռl+:�W�t���� ��c��C���U��h9��]�R\�T�n3�F�2��v�]�<'P��e���������>��m�Gdr˅� w@�z<���6��)b-��#�d�->� �ӑ`�d�-�T˘ H���,i�.̝�E�2E��)8�������5��=���r�s�-�>�ʞ�U����n<�GZ#�G�}ӡɂ��I�a圼L�W��cij]}���o�z}�^'Dp��"`�5K��vGw���������)N��z�+�P�� �8�O�\(8 �N~<yQ���:36{{�C#h6]���̄��^�����/��
���ȸ�8�C0�J৔����?g޴��:+����~R��Xz�N\"���CL>]P�~,��C��ͻ�V�<�� �m���"H"w���-��:k��Rqrp�좕�S��`8F�`-x�����j�K�bHU�;�rV����I^�N�vD��RO�z�:2-�h�]R�DB��>
;��"#���>7q�b2o�w���>N{���:Z1t����V�6���}��hJӱ��Ղ3��d ���,��<X�[�w9gu��[���j��	����U�n�vDG1�]�7��)��O���0�o���(��e侧����I�	��7�!j�eJ��u�u��ÖYe��g��v:`W���� -Jyv�+�H�%��J$�{�
�p���Vq�.H���U��7����2n���$�Dv�+c%��ZHn�J��O�8X@$��������d�����U'	1�����RmҐ!7�k�s!0	ӟ�QO�zm���W��8h�=%O��N�^"��C+h��S�ة�
0q �N����S:��v���cF��6f6zG����&=-ȟ'�<|B��j��˄��v���;B�8�� �4���w�W*���x���Ĳ�^��o�u�%܄:>����<s����=�����a�e��}g�DL�sy%��!҉���x��?��(B[d `ڸ�-C����[��յ��:��Aΰx���D���e�6������T�uja�,�7���j8�B�ԯDk�PVs��cK�h/۸�
{Om@��6bAƑ�����bX����R��L�v�8T9�$�s@����7�
�=2��F��=7�R�<8/�oGܨ�����(d��__�(]��c�-EԌƮ��,�_��}�Y>�Ĩ�ږm�v�v�������,�p����(?ȑ	��r1L��Cpi4�����{�?G�w:�'�L��&+!W�l%=�S��x�	B�x72K+,��Ժ�+�86Ӣz4
54���D&+��<��T.��� �9��y:��r*B�<���OO�(X�7�M;V�Q��|��K̹G���AW@��{K`v�hS�K�ؠ�`��&��J	?�hF�$MA�!���JZ
T��B��#�`��\�N+���C��xԷ9�45Os�k�Jǜ���AGDE���-+n����j�'��4ߍ'@����W��y4�������Z@��%&!��¶IQ,ϳ����J5��x)Ǐ��w"����jS��;��DI"4��S�HJ��`�ϝ���z��mǽmy�kp��Z�m��%���a�������9>�5��&�riS�-����?�+L��m���+�9���:��]��N@�o�'��,�R��Pn�ڭ���>=��?��v(ǒ7J��d���pO>ٗ�/&3�����慌�W&���g~�ӊL� (7�'����:��y4�j���SO�nhaBC94�:�6�ߦ~v��`l�Y���6n�qލL���>fl�"�x��٨d�R�8���d�\� ���N;;&�
�3����!_����K����s�גb`�#Z)�&�eu���g�ºق=b��u�����1�q�]=.�=lWRt?�s{��r%NS� c����#=C*5��݁��5o\W��3��qӏ��� ��O7�ȇ!��$j�|N�a7|Ґ������}O������?<fv�ҍW���,����m~e�.B�V1��ñ�����볕l�H�5�e�ݤʞ#E��j�!1�|'b�O��;Y�ruY@;�� ����?�����L$+�*gu]�)�������ě�����2�':���ؗҰ�}��&HlS����m����˞����޳�������l����J�D;�Or!	L�X�����1)���0	�r�ӧ�f������9����=�&��xed��3�Ŭ��;�j-Y�KG��嘍-��^�HP��u��Ȕ7(g�:�k[�!sL�!��2��0�/�U��qע�p�Q�~�Mlg_ʰ6�7]��ѯ�!lU�$��θ�H��:7(�wzۼ�F
z@�¤��x�z����g��l0�툗
�sa/QG�j�\Y��������]��0@ٺ&0������w�)���Mم�~$�bv��V���s�?<�b��<�iT��c�� ����4 �=X�C�86�:�|C� �*��ۊ��*�-]��k���3��q�D)e:�-����t��^�B5S�qH�4@��\$��}8�-���b�fQ�B^o1��)�Y�P�!�H�'�vMs�0���BXf_;����(AH�CAc�kHC��rͦyV�TTK(bq <KCy%Nhe��@����s'8�vT�o��1m���p:�Ǐ��P1�œx��L?�?*n��۪� �k�J^��*����˱�� ˜U�.�c�{���W�M��=
b����$h �Jd�M�X>��u��/?��4�vR�\�CY9ր9AE�Gvb��߫���.��08YB=���?��)��!���i�f{w��q͹��� �]n�m��n��jg��:M/�f�9�I	4��<�8b�Q�K�nc�4h�"V����L���ԩ�Xi&�qX 9F�q��"e&?�� i[�T��O�l���&��O1��S�֜}N.��92WCz�"�&�E�(	Yv�E ��.*�}̙�&��ᙯ��c�
��)XM���hk�oRI-e��	��H��`�ᯓ���C�
xkDe�#��3�����	���S*��󲲫�_�S��� �욼�	��!m����
k'�I�q��z8�OWZ�p+r�Ǧ�X���*�CJp��c2C�e�Fx{m�ZN�ͽ��-1V5�5�@���z6�)�<nB����'���G�?%��U��xG�!��'ѣH�Ĳ�x�|�Msk�Y�&+S�����NӢ;۪�c<v��n�E����W����N�ϸ�9�EE�d�xl���� ��J5ٚo:	`�4x7�X��É��Q��O�ĳ����=��(�mS���b������>Ba�R�0T�2>5��K��O�/��ˬ�']X��ÿ���4�Ȋɜnr�E#�It^��K!�k7�4���8.�gv�Ū�{�H)rB����U��|J�"JH���1D�d�2��7���q+;��X��V��������7_z*�*��x�XS�e�(�pDX�(!�O�o�;�x>��]N���� �����pFCZ�B��)�![dC0[���x]ׁ����$��Z�kT�
W� zׄ��g+0�"���v�Q�1�f6�u��L�L{�Wt�RSQ���t�?-P�z�{.8޳����5D���G���9�[���$xYk��PZ蕱��L܈$�)������g������E�@�OBY�J�	�2��<dV�=w)���9�Pz��h�V�A~� �����NX�`��&^��8�[~������/le��w���;�m8�%m^��W�گ�)	.��������!$��O�A�@]ٻ)�[s�&Ahӡ\&�X,H'�Q9��YV�*�I����6�q�����^��9����Qb�L��Y:E9�Px��s��"B/�|��0���v�f�O����C����h� ��W��O�T�}&I1��'��O����u%��lQ%�Z)�U^��6/���9��B�؜���6?F�]�����H<����Qv+���^.�>���ܗ��/���, J5��\�c�a�4}�w�מM2)J�g���F\T�Jd��哰�ݹr��zԕ8;ga�6��c+�_�!��>��ګyPV�N�}�.�5IU4Jr�A:�1a
?�x��Ox����@�;k��������)���A��l�>�����ѷ���,J�%�a�\q���m��]�̥"TyX�e����7�S�����0�ן��v�Os�
c�"���z��6�[.Z