��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D����gP�������������44��Pg��w�k�n�L�t�=�ʠ̲J�=�	�$tG�讧��p,��sC��Xu�_ S�	��mZK�qnu�*u"ǋ<�L*�2S���!��i�އh���
������)�=k��l��hx��I��} ���l��CaoK^G����F�HE���}�-���8���C��)�6v��q+���BɃ״��0�Ўl���Ax�`93Di�j�]��0x��uHo8ȁ�h�+���]�,L��uS��|�>5��9�8>�U̒ �|�o=���{�
'�[	��ԄgI.��Rs���Z�GݲB�_/h�_g�ˢGmYAa/E���,Ӥ`�΁b�d�@��+
��kz<ˤ(�w����0C݊��L87�C��������z��H�w��ڻJ�:>A��>I�B	�KW�-H��
 �ѶJ��;�\�16Ji�,�z}�:d�9E��_����Z���o-�[Ɯ��F$v�KG�%Z�:�oA4w�)[����:��z�X�o=B�e|�_2��ͰUSo����I#ظu��#x	oC}�v�%����KBU�2 p3 e�+�0ʝ��l�;$랉�A��t�h�?\�<��d"]���xuB�@3�{��e40/���GC��������ھΛ�HWR4��M�q��q��x�Gf�5�AW@{�-��LX�d��փ��Z�$�|�t��u�z(t�]7C�ua�Q�t��>l̘�9qaD���5:Ee��LsQ���荌'�^�� �̓�4��QɊ���	�<�P���yJ1 7���x-��2�.�,�Z,꡷8 /�{�{���*ٟw�a���r;T�>du�3����$}����~E|2�E���'Z[�O�sA�����$�W(4�:G��Zq�! �F܎���i-���_�b�F�ʉ��"�5����TN0�����,�����i��SR�>��H�nX��cA�<E��RF�k`b�`N-˓S����G\�1�5�s�"D��tD�6����L
�������v���bM/�<��˛+ts�`Ԙ}�|�l\�d��g�|���tm��8Dy]�s�ƒ=yl$�U�9k�rF�	��:��<������MuC�����C�WbNḐ�S��?� C˙I�Ep�x&۱g١�	�w�s���[��3� 
��E�a�{A{Ae�#^R�^(�;�q���(�������J�S�bBo˲y '0^.򩶙-w%�π��k�i҉��2��]ԟ�Jx��++�O�����s�M������\�sG�w�s����#m\�{k�Wv��β $9�/��Xba @��(Q^��Q�Y=:A��',;]�ų�M9y��
�a*G�yy��}��eҦ�C�9k�a���\u�?Z�e'�h0t�����KR�M^�٪�2g0<{�[��W8o�$E:Մ��q�zqU�I�l
.\�*"\)h��t^z�6E��]X���������0+L�t&Bc���m�d�&;6��}������!��pB:E!&���7�t���7��Ǡ�"��ݚ�NDjH"���Yl�0*&�G��|[)|�%�����r�4��ڤ����H詼HՓ^�P�^�h��A&��5��O�=�y�?&�r�O�8a"W�ˀ�F;W�ڀl���yQb:�f�.��w�\U�ʬ��O�p���m��%=�[Y�����5FqI����b�L{r�}6�#>JK� #sr�9��	� ��T�Აr�&����3}0�l�\?���m�vR!!mN�� �˒���u��P1Xk�=&'��q�E��m.�{9�*�Fne���9��Y)OM����*b�㷍$ 료kl)^a��)���
)��r��h�6�,-L#h[��mHa��-�����������"X���F��.@�U�m�L�V�`�ʎ:[Lܧ}������X�����s�r*ߴ��&�Y��ԬϚ?Yq��2����x��_��nOsJ�U`�2����rh�%��a߻�f� �%WD�.���Lc>]�z�<pd? �Z��O�ͳ&n��=�N��-.�)���:�Ïs9�7aя�\"��j��I��O+�Y�l�ΰ�Ol�9cl�$��߱"�	���T��on`��~[�Ù{�0:�t���!�<A�rх��x�[���t�5�;�q�+�����E��%��W0��F�rfF�_u���tH�\h�G�_>&�S-�Vօ���,��Jʠm\��|*����?o�rY����V����S����yT A�,�$HF
�R�[������V,^6�v��dQ��Ʃ�6�X�bK��
���m(U'�y|Bţ�*%}.Ao���"�%`�V��MerV�<���\�M�:��c�{4��arr�5U�bqz�=���-�a��ї[��e�A��$�uK��XJL�cfV���/>W��kL8�MH�fβ��v%@��j�[�>v�Y|)�^�͇Ҧ��W2��۞v �f�c�Zs�B/A�_�Z@�_Q�`��p����e���$F�XA-f���R-���MW�»f������Z��G�"�q����rab�)�X�5B��q�[C8��/����i�̞[~7Ն��v!}���Z�x�-s�mZ�lt�Hb���U�1�zZKn�;r�
P�8U�J���h��멛�nV��p�d�>u��X�6G���u��H̷��3(&º2���O��l^�����*�A'r-��{����1�Y2Snq�K��{�Q2ڏyU��g�灔���7���i��
����Y������{���`�A_`�t�OI���c̎���B��0