��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�Tں~�ImW�.�^�ᆹ��������]��%�wx����xeՍ�ϡ�&JLc7e��~�'[�b(�Z��M%기_��H�K%_N�kV�.���a�����F����B�u�E�[�D��*{2<(ڡ�KiNO|^'�`�Ơ1Oh��i��=4W)GS���A��+�O����x��g"X �Ӫ{T�E�T�G2	0 ���F�h��E�L�W��Y,N7b�!Ů��N;?3!�o��Y"�@�V�+y1Z���Q�E�H�+�U+�ϛ8k�!
p�A!�	'�E�.F�~��]x��:r�i��J��߇B�n-g��>ڶFW�XX+_YfS�k�s}�,�rR
*�����=�N��#E`M�0�8f�d�2���ju6<yC��Q*��Љ�/�Vp�� `�ܔ�e/3��&���"o��'\�Yb��
�xCy�v�1�n7Z�_��i��)U�)>�>C�ϒ������a;*�-��-J�`Z���S�� �|_lIi�ʼT@��#8k$F�B�����
�@�� ;��g'�n��U���yƉ �n����7��0�p:����;a��}e��;�1��::��Ǜ���%�x�j�@6h�Pu�ԳՕ0nf���gkZ;�����>�̲$�M�,師�!vlG��i�̰u����Ⱦwɨ�S20�,�_}F{�s1���+������а�pU�W&�>��M;��*���i@�)��m�\h����D��+���{����i�b�y\M�-6|]�dv��N�vX!���f;�i�`�)Cx7P$��;��T^��]לO�oZ����&�22°�,�ysk"�R��L
"���e�>����� ��1�v�m���)�(``#�R#OVif�9��f���vfƼy�f����镆Js���ƞ{9&֎r=X�	�&ǔ��A��:�O��G鍄�&����� ��u;��$"*Jd���3�*�����8�D$�t�p*k�@�����3�DMB���D��f6��U".�km,X�y�vC(��;�4�.ֆ'��<���Ր!4U]��_�3�j-�D�6��������̏t,(Hk�5���!%d)x�����n����J���u��2흧J�K����%��LQ����e��b��_>2�����&*z���7L�ʚ��a]�����.�����a�����y���rN���r�"B�'�) ��u�#�I���/�� x�Α��Y�)PfUB �8����F�N~�+��Yp�`�G�g#��'��}Q�����)Mjy|�?^��t�q��{`��O*'0Ĳ1�j�R 穞�S�U�X�lZ�>�kj_���o�����z�gg���ƾ���݌h�������ɩ
v�i�.2��?�c.E`���d��&�eO"q�b���$�܁�n�������H�H��|q2����Q��~���������u�k�Q�aJ'
��|�4pɏ��� �%�D��
�NO������MYB�A��n����h���'aȿ�� ٻ9E�wu� �C��9���m�yղn_y���2#���e6�E�ʠ�����ܛ<�	�=PH�W��A��]���Qݬ�vW�&y>��S ���Z�J�a�^u��(�8c����j����%F����:8m�����q��fa�?��|%�]ƭ�$���S��J*�=x��~:(h��{ad=��?պή{==�� ��t.��g���'�;���c���"�\�޶�Xg���Bv���m�Pg�I���q���Wd��{:�m���K�@H�<W� +����;�K��fH����zS��ʲ�Brj��G��{�~�O��he�b�A��@,y��Ejk�Ĥ˧E؍
b�[��(�3�e�m�	�Ѓ��ȩ��#'�)���S3�w��U4��s�듮랃,��K���Xf0�|�=xڬ���v���=T$�8�c"0ԕfG��:J݉��fZ��H<�w���a�C��� ����Om؍��Ø��2�L��z�Tr\�OV+���Ɲ%��ҢŜ+67_؎;�G�a\��u�Pt�  ��t?ܱ���-pzR�Z��~#�!��'�~n^�w	U�G��;����El��%!*h���
�`�H�^�#s��������q�.k��:�vb���,�d<Z�(qL�������K�)���hC��gk�6<��gX���\R��Ϳ��.��h�۽;�5����|���|��O\��}{E�������&�yߴF���>#�����f�狭(k^�?�!e�L ć��!��PԦrk��,z�"l�UN�q� ް鼼?��ԗ�+Q��l��ū�0䟐��e0�[T����aܓ�F�Oh�c���()z&����e/�,�8ئ^=ؖ~��}iy�Zf�+K
����NʤOo�	|�=�6ă�8��#�ͥ�B�R!�/.,TG�\����@�<�÷�;Ui��9���c�؞���ϗ��Y��fTW=�X�OC�0h�}kQR���A�{�N�)� ��<�M�U��H���Ú8�)�M�tvʽ��^�
�5π�tw�7���)��
��͏���w�_���Gv��Gc�f=R��c�B�
�I^*��l.��R����,t�&o�/�1���8�/��Q$5��i�dp2�1^�§3w�ʌ��-*Awg��u�1x�Xr�	vB`^w) ���D���6�4���B�J�u�����Ba��_O�+v��;��"��貋^��v��$q�뺷4�&��S��y�����1�8�m>1P�@o��ͳ��|@ <�(�.����л�����+�����6�PG&�����o�����?���&�TM��	b�r5�K�W��W! ���&S��RN�4V�����G�M̈́�}1�vIP��qE~R���D����4<cE�}T�7��Ǹ��涠x+�՗,ܹ�ZɺZBM��6O�N�|��4#�L����p�&v���ܹ��Q�|d���g\�,��A},>����w���?�=f(+҄�۟��B}��̕߁���������z1�1�0�mn�����M;n^��Hl�V�Q@��[�<ʽ7�KF�X�M�fG`$j�(18�`���Oc�8ō�t�=�����ж ��0:E^HE:���$�s�}�0x�ɺ���d_qu°�4���^��J�4��=�'���^M����s�S���*��s�Xu�7��d�/f�����F��ԯ�U�"�G� �%�|[o%�5U�\ۉ��W���y" �!���Ѧ0�U��1���<���a� �s~��cE�:�|-�G/{OM���:4Eϟ_6�J{4��j'�t�q�������c[S1�n�i�,t��htΚ�Z�Tw\h�YĬ�"��9}�z0����n�( K�L���hk��D_̍Y��tPu%
�[^��e�ҋTrg��jà�g��,����Uz����x�����=��x-75#����v��B�٩)N��@Q�\���,�?�^O����c�����
f�ٕ��u�֕E5��ꣾm��}��C��s�r��4,�rԶ�ͨ�S� �&�bI��B$�U�֋V�dϟ�$�x����~?��foi���������d��a{FU��<n�C��m�~�,Hu��8�C#�P,,�/�_���1�깘��3�� ��- p�	�7`ћD��s�9<(��ބ;�����9��`e��:�!F�2?UM�� b�#��VFuU�+H�����:��?���}�ע�+��è&��blaL��}d#a��`��^��t+� ���I��ݐ�ӣt�lS�TKz�t�h@���4S�c~`�vG�qW-ٕnFX큘_���e9���ք�	�*�[�Bid�kJ����-0�w�����0g}�&,�Đ�@�G4l���G�>��r�%k�[��Q�u.�l���U�]�=�5�?oq`��1�L����Ն���sX�/(�:N��ҡ�L$3�c�(�r���wRU>��[�c�f���6�R��1W� YPP����6蟭�LE�]D�oXk�V�|�9�R͕��
�f��]��F{����_<����˘�^�x�Сb������I���gi�Y�j|r���LL�m��6�NzW@��#�$9�ӫ�����b��Y�%����iG��ǀ�CD�俗�	�R$bMh=n'QX��������[���tR�<�w�;̛嚨?�i�����(��������0�)°K�B����M��m=�\��A~�΃\��FGtnZ�nz�Y
by���+������X�#��$`LCL1��B�&ALj�+O���hȵ�i��/�U��P�%k�˗ض���t��HuX��E��vm��2
/W#���RJ�7"4@mK�g-�i�˚i��@�qr�����7d3ɦ"l�C�h��Ӥ"�a@�~Y���naD=�J6�R>j��g�G�+��/Vi������*�z��I7�O�������<����Q*�Bi�5�=�z9�h������#f��U.F �����4w���p#��J�z�dw��SpdN\x�[�p���S�JE��$R�K�U�S�]F�8�7dlK̶5ctl��&Ol��q
qG7L�KT_�q�� J���Q��9�@J���}2�{��"���b���z�b��`�c]h9lPX�A�)����y���c�4��ن�y�7�YO)��DyG,?���*�L�#'�hګ˶*���h]~�kR$�fx9�?��yS�<�,�M�9�������y�&���0�r�M����Ʈ�(�����0�])��k"ԖK�-�����o�ʒ<�̠`�0-��YOB$;N~Ԝ�W����"ߞ�so�Z��L:6�smm���u�m�����iJ�{+�^�L@�,0���z�ZE�\�Ep�V���[GW��%�ծ���ȾF/��o5ґ�W��T�FnR�A�`m@��ױ���f<�Vm��,���`�`�j3�F���U(${��)��xu�8#7w<��j��4�52����O)J���x�Q_�DW��m�e���gTP����a�P�(�DiPC�o:c��7��B�?�wYW~�	�_�Mv�B-�F^%����r�2���3�&�ER���R�=)���h�V�[�V��չ�z}�8�H��d�c��z�;G�!`/��2?�W�DkY���R�X�\��y�{s��X�'s�)p
���3|�^�ɆR�ұ|gdP�j�����@v��5X&JS�ユ)��Yt�X�9R�#"�4���6��r�����+u�@T3ܣ��nf�x�#���|��,a��>��\���D���0ˋ˛i1���}��1˳ 'U|�o� �-��1�W���	����kh���3L܈3fɣn��u��娫�͐�7׿�%�]��֕#2.r'��5�Oٞb��?bE��I��;~�6�+�����'~!Z��+ʜ8#�`��9��V��ϯ'11��D�O<�/�-�=���Jv6b�QfE�\����R����<Ȑ��{Y�{���,G��k���!�|T��ǃf͓e�CK_��21!��*C�������7Wu�fr�s>Y���ju�+]:�A1� ��l'�ad2/5}�b�tm`Gs���׉�a�.)uѻp7=��h롕M���-��oM���^o��?nk�G�?���?զi������)�X dⱧ	��a�.��ΚvX���ɗ��%�����t�2�`������z��;�اз���pe����?��}�����g :�k'�mஆR���焽������N%�2����9��D�O��F-���\;=bG <J7n�FfN��=�j���y	:�G� ��s��U�L� گ�S��Ț+��d�mJ���4Ws�f�Ot����j�Ń,�ȟ#S�=M/C��� �������[���M�����₌ԫZ"PW�!�Xd�N���*�T��� 9�r[RC|��M�n^ց���AXꭓ"ώ0�Ǻ��_drG�"�`n��?B	�#�v��^-�Y��S��'a����ҕ�=��"R��;��=ë�-&ד����I������З,%�PN�8��K�;}���'�o��c�P�4�6K������M?�,��o�O�02�&��ߎ68�v���p�o��A?pc^υ����o�8r^d?�Su�u�����A{�f�p��,����z0B/ܜk-�ၝM�6�4wW��q!"���V��\��^��ǉ�myĥ��dm'�'�G���őM�A)��%���V$*�Aaj�P� �,H#�����R��V�ގLb7ݣ~3�Hȹ����F��;�*_�Ra��W�\��P�CW0~:��?�_��r���h���/'��bto�>�	-!�D�_�O)ڻ��Yv.��-�k/�yv������ob��t��z��D��--�񌊌�@�	R�=o�?��}� HV�;��l�E5y[�� ����
ڊ��o���WB_������9�ڇ)5�Z<��g���J�TP