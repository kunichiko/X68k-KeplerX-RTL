��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D����gP�������������44��Pg��w�k�n�L�t�=�ʠ̲J�=�	�$tG�讧��p,��sC��Xu�_ S�	��mZK�qnu�*u"ǋ<�L*�2S���!��i�އh���
������)�=k��l��hx��I��} ���l��CaoK^G����F�HE���}�-���8���C��)�6v��q+���BɃ״��0�Ўl���Ax�`93Di�j�]��0x��uHo8ȁ�h�+���]�,L��uS��|�>5��9�8>�U̒ �|�o=���{�
'�[	��ԄgI.��Rs���Z�GݲB�_/h�_g�ˢGmYAa/E���,Ӥ`�΁b�d�@��+
��kz<ˤ(�w����0C݊��L87�C��������z��H�w��ڻJ�:>A��>I�B	�KW�-H��
 �ѶJ��;�\�16Ji�,�z}�:d�9E��_����Z���o-�[Ɯ��F$v�KG�%Z�:�oA4w�)[����:��z�X�o=B�e|�_2��ͰUSo����I#ظu��#x	oC}�v�%����KBU�2 p3 e�+�0ʝ��l�;$랉�A��t�h�?\�<��d"]���xuB�@3�{��e40/���GC��������ھΛ�HWR4��M�q��q��x�Gf�5�AW@{�-��LX�d��փ��Z�$�|�t��u�z(t�]7C�ua�Q�t��>l̘�9qaD���5:Ee��LsQ�����yEE����%Zg��Z�؋�����_Z��JC�z�
�T��%)��G�_mu=_��w����M��\O��lw(z����tВ�"�׼���E��ς�A�qy�<����1�˹[��W�|��Zy�=q����H�������t��y����8�̈́�����<u��b`���lcH��T<*wi��OK��i76ao�3��+�e��i�M��NL���S�p���۲\���-�@T�WKC%�v�����(�ȯ��#̴�ɦ��ʫ�����l	��H��6��k�Q�i]�8�.9��8AJg{�g�mwP����Dt�X\e·��h	i�]S������,b�:2�p��'�U���Ы�	������Ӣ�qw��jU�k��,B� 8�{��G?Φ�FKj�&�������Ƽ3u<&H�P?���ٞ�AOgE���<Ѓ/�N�7�Z{<Bs��h���q޴�QԿ]͗A2��0���H��%Lp�3�
 ���=+����'�!Ν���/ �P�q��Ы~s%����1�q����������Xr��/�������Ja��]�Y<���6�D�ź�<j�m�4k�d�YƆc��WFث�O�er�l�Ve���1��~�{^Y�*kZ|�D�g�Ǡ��M4�#D+�g���N�+g��^�u�l�i��$�O����msL�E)����I!����6��S$��E�5Z��Um�XMz��>?`L�&�QR�����Oa�� �C��w�����aH&�eY� �jm�bW�9���(x��������F��
� �c�u��r�;��Az������e�nZ�GI7�6�@�y�8��:�@'� �83K�cK�p)��䆐�T��#�&��6X�����B���5���������Zxw(KC:�U���*�Ryk^��?Jc��5��H��M���M�谷������$zr�H���	�H���`����zvLx��d:���@��y�T9b�8T4���|��tO�\�y1�
�������λ���<P&�)��U�T}M�-%��N�S��nt�$.�l���\�3�f�Z�<��U�)p��Q��ŮJd��H�<7��z�3H,��c� ��-.g'����Qjj\S2���J�����	)�l��aRF����g`W���g��h$��ٳ֦n����/(y�T���O1ϖ���]���v�9�\�iZ�Q��)+C��`�g�Ӫ����i�u�D[&��{R�[t�أT�|�A�X�V�m��8��+e[_�|M��9^��3�aq-ї$�����el����� �����vQ��?(�W�^�D�F��",�N�h���N�-���<�����H����r,=d5�	�d�	|�����p����7�1��2����'m3y���P=4�"l�9�����/���n��者ۧ�t(��>�E��������"C�w>�m%��OJM?/w�#+��⨪`ƾ�tJ>��_eM��u����#�k3���R��]�#J=|��r׆��u�md=�bv�n�H�3�Z�sR�H����"�+��{��dC\�7x��'28�������3����{W
��-�3�@$R��-�x9�V�N�a5v��$,����}� m�×X�P�-�ћ=�q��ZY�m=���p�X��-�	Q�O��hkQZ�U�XͿ����yC�2�ƅ��i�>?rn�P�CV�Fs>�!"��!���5Ԣ|Ps����3S��TT�/?�6�̩Mp�O[V�o��gx���#��Ov~�KS�r��;�N��e;��Mp����N�ګ ���#��PX��A�8�;p0����3i�4�p�ھy����p�'S��#�������q�^b`%�l�I^ˁ��W�$*v;�	t��6[@c���d���T͑������*H0K?���x|��d�mt8��ȟ�l����KAb��rl�r40�B.H����~�Hf+j0<��E�K�n�3����Wn�i)�dɰ⬴@�#EBv�p 4{����W;�+�m%��C82��h��w�A�ih���OT�+K " bs��"_�DQ�]���b�V��[FL�/��^c��&���0�+��k�W#gK�fɕ�j�%c�]����#)�#Ut����.O��w��u���$~�y2��ع+�d�M�|V��4s�IܹL���%����f�R�B�ڧ�5�)�r��kkH�/�kLwS����q��{��?��v^�떩�/�C+x0����5����Y����҇Y�8��-��,�Jm�)m�T�
Ga�4K&;�} �7�KJ���րx[�^�5���y����之�sGl �k@p�k��n9g��ޤq�^䇠XԚ�ݑd�PDq��%O��O�]���w3i�w.%4��Tu\\�וn��� �y#�HRJ�̿�?���wacY�=u��o�L]�G�b�fy
z�wm�w��~�g�����d�s���4��_�'�6 w�#F`�g�4[@e��r���8����h<o���@�6������h�+颋r���8G�X��@��h1��.d�&��>�+CG�H/�((���t6��"k3Z�.��1_�Ӓp@�4�T;�\����
{���B���v+(�^�%=�A�s.8Q���WxԎ�	�w1`X��Ť�����C��nV�;T�I�mҠE��k���k��N�el�.�	��sd�1s㍝�
���h&�m�ar��NBOT�|���R@�>��%�5:��AX($]��m�[9B��!U֣'��t1lE�Á˕/	3�%yF��3�2�L`zw�p��E�f�Ya�![9:%��e{Ԣ��%�����]�[�F����_�\���s��8:��K䨚�#�l%�\��R�����\��ۢQ��]��$!�fB�F��8�d���,�����.t��9_�6���m}غc�pc**�GJ�{��}���*��"Ƽ�YK���v����V.:5����{���7���%�k5y-��
�$��Ъr������!�%��4HY�}__4@<�NEm܁�B�X
ў�ߴݟ�/�sI�b(G/��8/���D��i�{QG1.�ؘL�{Ig�ي��;£�2f���a�D�\}\om-P��~`��֫'2�WS[�*�����9`D���ˣ�Q�ښDˉ����҇��Z�*7ա�x��Jq�/�V�]D��*{+-�?
��6�Hے�=�5G�������c�;BY���2��z��{�b������������	׭X�N����̅�%����PLc��R�݀O]�� �@O�0�b3��k��͛��cp�x�U�%�R���p��1�3���ߌ	q}C�tfL3��Xd���D�3`�J �F�
;��!���n/�yg����dY0D��w�E�V��$O9FBHʠ��d�>j����~D�@�.�a�����.�(�O/�S���T�IĎ�dPLeoԘ�۩�9)��mF�j�n�uU�x��y0p�*�(����U�Q
<X�Lz�����e�(�.��Ȩ�J�̆���Ͳ�`Г��=prjH�-f��+XВ�	��=k���A�u�ut1�ږY�W�]Y��
�����r���%ҫ��4�\� ;S�����<�G
@̀0l�Dxg`���"�y�xh�Ispn���"H���ʽ�@�A#��J� �n�ɰ?4�eQ�;�Ds��8�/�TP}W=��$TP�]BW;@�d��g�(u=q}>�.fX����E�Oe`mѪjl3n^]�1S����!s+7I���>\Ǝ&%RS�?;aS��,y�/��^4/ׇuO�\5[�� �$u��`��,p����ReOm�q>K��nKM�$U�$���ʑ��M$J�e�$o��b��鵟"����p�䠐�ue�}��l.h'3"A�	�)�Ȝe�U���By�rV��Ϫ�^8/\�A�v\׶x�
;���f�>�KP#="M@3�c_�����d��4�|by�.�w:G�E�9�i���4��r�P�s}�K&�Dښ,	}��vSCE:/"}$'�e������_��^׶���@���h��"��g`��9�
Km��/Tي���g�����u�:�*������0�9%˙�o�������rh���E4k	s�{�"lm{��|c�U��\��%a3<�Y]�L����l�%Y�|���+�!��G����)EbӾvQ�3T%!��pݜ]VD���2߶Iv�z61{�i�ƺ�������kt������č�[\����|)y�%��n+�^���u���	�������s��h�~��eмG麽�!{�k�т�i����X�g�Q�@��W�?=`����cJ[c��r�%,m��Lǿ�ݰ�	�8&���H��_�=�a�����%$��������/N�dN�ل)9��b70&��V�X}�{;T�1���P�"�� �&�,^��U�� e�R4�r�*���:R�MRʰ���I]�ybӚ�[EH0�5«��^<(���!j�-ܰU�~��F ��K���U�/J�wPv�� ji�5y8�	�1�i�b���D���pFb�uA_+�cfD�w�ӝ�ʆ"�r��u�S�@ǯZ��_,��Hʏ��1F��Ҭ�����,���������7o� ݭ�s�S,f1F��,�-�U$�Їܱ��>�<��c�Ȓ��媌���3L,��oN�l�.����r��ψ���B��n�(k�q'�d����"�ʻ��/��\�@z���F]��Cڵ9l-�z��n�c�=���n��s��S����|�h�5�%�-c�� ѡC.��y��N�ЄE��_�ưc'i�!&��	p���R�*�՘�Qې�|�h*�4p|"a![,Ӝ�t��-��k����CHvR�Q�2���V���	��؈b	x٣vp�E0��)�
��?�l�i0W�X�����X,O������")�L����d�Gr+503������Q�+��-���(�i�")a_e��]ks�3/+������n-�aM�O_?��1�A��Q�*�*.��r)�r���̟|��bċ1�d#�j:�B𣮫��q�C��$80[���X&���$�2|#W�F_ 34�� ���O�1��D~ `}�������4x���X���xn�\
l��6/�A�=���K�m�?#;q !O�Al�u����}}� Q��E��T_��(��M{�yx���N���<*h��毝VD�wm�Eq�(��JJ�eT��}�Y�Do�������Ѻ�	D���i��,�N�5��Z;��V����]�ÑL劑؄���ǂeH"���{kU���s�w$ި�������s�Q�P�ش��Ū�.caB�z����Hd6$.���Ω����*�kD�a�_�4~�G��u��T)��zY���PE�$�Gb�ez«�� ��G�Sfc;���+��1����&�S����l|tF��9����$ۧ9�*��9�qp.Y�����Z4�Vy�I��h���!Xv����g�g:LK֓��J��]M*�&+n��\�n���[�7?�5�nvo��k���TC@i�oz�����TZ.�p+���Kƻ��sL" A�_�������|ԕ]t��C��!�}��-��d�B��BA$���VCs�-�N	�S�oW�/%�j�&ݯ"����QE�\��򬼫���%�!�")�jnF?��0��IR�"8���*w�S��D���fuCW�u-h`X�li|ȭ���?#�!,I�U������:�Q-Q��I�}g���� �y�BvD�����U׉���h��j^���������1��o6S8\��񄫯[�UN]�IQ�tl�FK�|��������ݠ�rI^0�rU5���[wpY��?gd�����M-1�O�س펴����#]�c� 8l�4ɟ zv��jsF��y@���W^? ���z���#��Ǘ�<a���55=�ň���~���JΨ1��<�3K�⻳6�Li���NxW�S�ť_��f���V�{Q��~= ���F�X&fv�G>1,o�̜e�T��?m��|��q�n�����_�!|	�+M7P7�V���r��.N�[
k�:�����RA��"�W9B#�Vh4�G#�f�s(Bf�#�#�K��w�s�:���O�|���xh��[��c�n�p��/��tMR6�V>_�>�����'��	�@�*�4m}$1<ƙ��o��yz�|�VUYĪ�k�9
��S�^�}x���x�-�-9�����J�����d0�X�D�u@��z�Lp@��AS�'	Q�S�/^���x��V�@��>�]���|V�o���Ta�Q�|mD�PC�nzt��/+t�10�f�l���5�ǎ:>$��B��gC߹�����R���w)4����i�34���#
��yN�9U�3��a������8�;<�u\� �1��Mn�eAE�؃�r���-'R�t=C���2�5��� ��e�nLj<��u��:�9�P`���&���݌��5 ����pOLO����P2��`TcVhD���I�Lp�@-| e�f�=8�z@����٫[[�4=*b�A�{
l��
�!1e����ˆ]<:�zv���q9��`�^�+X�}�j�#M�ŀm]��,�Y�"mɆ��m\~�or�q0����^ް,ϼ�=��|A��'���2(���j�ǳ���9=_���r&�痸r���,+-黠w�l1n-[�����e�̄��n�U��D��S����������w���_��p�6�>h2ȶ�ڃ+{��������!4��AL�7���5�v��K�ù�F���Y��V�;��PNm���c�[�͋����%��{]WdEE*���twja�@!�~���7_f>m���	wo�V����H0�V�F`_T1��5+�<]T��L�G�|iP�]��Q��G�Y���e�d���e�Y��U�d�^%���.ʜ yE(�I<�6dr���Íٹ'��%*�BHԐ���C��u�<�n�8 �ob���:�p\疖E�E�
�o�&�/({�D��œ�W��M��֕\�iP�M���0B�)pGu�QZ9D�yq���`n�-��j�k�t����؀��Џ��4��xÇw���I�e^�� ��?B��Qw;����[BŖ=s�X�5�kA�zs �%�h`��R��,�w]����\z@]��\"Rv�ԕJ8�_Dn�<���x����`ɦ���9nۺ�E�֘��]�LrK(-q�ş��R�6��c�pb1���B���^�Z�q~��o.0�Ӆ]�8��:���p���ON�?ζ�=�����t��]Ӣh�e`�
��%ӟ��sg(m�NN� F����QU����o�g�oU�K�"�hA`]+�#�
�/�u��N<� \vz�c�����r�� Յ�LM����R{E��Z�OnԼ��0DXBXIU��5������g��4'k&����I{ߏb"�Md[@mpFR4�������{�q#9J���GB����񞧥/�z�Q���7y߾�zB�������x+�5ǧ�%�Vؚ�E�A_T����J���^v�y�=�&�z��T�t0�}�?u����َ���S�yOs9Ŗ��>��O���Cw��	����t��G��u������U_�:#��g*A��ܤ�W�0o' �1�[Q8������nx���WQX�u�û:,�?o*´�*�
&c-�.�o\>l�1¦�r��TF?�;[w�6�XPme,������;���Ꞓw��k�a�5��������,�L���輍�� +e�q��r�AƗ*H�n�s�BO�|eϰK��D�6�t���<G�d���|�U�3\������D<	Բ8�2�����D�������.�q��2������4�A �]ҵ��V�{�A�4���/���T�f.ІB���gP��PFw^��P�@|_��+��!�h�Y=A�gS�|�bG�H��/\��f��r�m����=�$Y5�5�3���0�jbsɷ�O�z؞װm�Ƃ�v�m�'m)5W���� ᮣ��*�rX^΀݊[,���Z9��.(0+��[�cuYN �N/��Y�e��<J���K?\��x��T��YN�"�d?�Df#���Uq�			Pn�W�j�%�b�Cݏ�҄T��U�4����P���1�M��6F�xߠ�pV�`.��C�����$w�V���k2�ˁ|�Xv�~�ʧ�N�e�ܬR��� fS�x�����'�U�aI�q�I�2y�ɽ���9V�9f�L�Zm�B���]�K%S�y�I}��]�����d� �����+{F�ݒ_�/�8r�]:S����|w-�0AR]��r�?7ʪi�o�/a<���*x�U������JE5�|�ݏ�dmD�t�C�d�
��yUD�A�i$)ٱ_��R�b�Vڍ��6��>Af�v�U�C���K,��o��̧�r�T5��{	����:��=V�u*�v���z��6Z��n{C�Qͭ�p?W�	˵��UZ ���>U>���7wҘ�@� �/�	ƌb��p���c �u�ZE��M]����6��<���qUڜ��E�cߟ	T���G����;L7�1E|�J	�!��'Y��!�&��@�^@ �_�4֑�h��%<׍F�ʆ��	1�4��Z�<Y����=ކ��$-A�"h�y�A>f1@�8���t�K88��� ����$K]Њ�l1��o�0}D�ǝZ[Jo4�-L7)�x_>(Gm�8L�!./&7_>��f�ws�i���CHè*�98�I�*��R�S�`�S�]�J�'E�+C�R2�Q��_ !��1�Ŝʼ<�	5@�wj����r
�.�w���o�}����,��9��q�ݽ���@6eR��������A��5v�9\�7�[xd�)���?r�%���f�o*�l�r�p����y�z�/��(Iqh�:9R��x���Z;"YғX���wE�<b=�͛�?pGT�hd�E�.0dx�g����)D-!� ��������I���j_�N_6�#_ Y��q\�[�Z?S���D�D�ޚ����bo@��^�o��������{/��G��h�΁U��?�U�%��?C��!/�w�m�K����M�J�9���{�w��^��@:��s�I�0�S␰��h�i���@���H�`(�Wk�Q�ʿ���T̷������<�k�n*�&̧�J�.�d0k$~��J�N%eD���.� ���z5z긣&��L���`Uᣆ�`L��q.�dgN_�7�n���I�Eg�UQs��k:���@�u���FN�Q/�͈����c��*����_��w����S��]�n��ٖ��K���ɡ�7���g�{9�\�-`M��z	lk���D�VmF�[��$�m��C��*_�]E1�7�"���W�2t4�����$'ߙ@=�Y+����Ƞ^|�~̢f����\��5��X18ɹ�~>jJ���M;�yo�[\�=����|�+ �B,�r@�1\��@�N��D��n�[8e]辨kM�?m�.<k7��^l�v�t-i�!��Zbk��;���������L����v�}�HS R��̿QVqZ�;�M�&�ǐ%(���L0�b�'��ÔCz��3�F���
-��ה̉�P����Y�$�@
���/u;�����8�k�G,���Q�3~^�bo�y�@q&P_�7&7���W�5ibLd|���RDL��\(�B��.*c^�V�W3���_����X�].O<��E��x�B7rw:��H<��#���W��X?���+�9��wr��_���1w�c6m_>�R�)��e��2+ �H������O��m6]%З�dI/ޓس1O�H�?��5Z���l�u���(w">���H 4'�ь��Z��w��&��θ�
V�mO&�mگBӮ~)|32Uz�^�U��%�h�^�N(�@nR)�W :@H�k�:0E�`�-r;g����Z����-:5��T}'zB8$n�+�ظ@p���H5vR�J���?��gaK8gC��Ez&���AV�C�=�%��X�!��r������Ul<)im��{�Zm0:��	��^m����R5�d�3X.�qgT||�	�r���ᑚrv�!�y1 ��8X6�;�,�O�ڼ�v��4�[)���y,5�9����Ӽ�C�L}c?��:P�֖ELo�ң�S��O�KwH��t9�*�&�9��yh>�H:%�:&�˃A�I+$0j����*aWĢw�'�)�v��n״M�5�
V���[[�P���e�ˉ�hjU��JA����v�O��ˁ��>��d�����:�1����PGU�g�gx�\��:���^�Lpk9s�j�}x����3'�0y��xM������.{�N��:Z#�=�4�ѩJY� ��������f�jv��~|�R���2�97�o����,b�|�`40o�>�1���`�D9��+a�r.Ǫ������!\�ǈ4�d0�e�h��$��z�u�F�����";���!_��m��o"!%�����_x�\�m~��2U'�4��꣬��؜n� rE�@����g�p��<�F��-��Ӣ�n�zl�(�ٿ27��+�s	v�����2�w+τ��BFˀ�H�r���o���|���Ɯ�)��l�L_���U���o7yYo�n������C1qf�6��ǏX�R��)�>@z�$J��*
Z��lXc�d���P:��("��Ј2���0��1��wS��� N�!���#�.֔լę><�O�k��,�*��,V����W�����-tջ*C��&,�K�d��) � f�b���R��+;	����Z@p�ɝ��i�
u�z��n��f���Ba��I.��C��[]v'#3dWlS�l��~��pgm㪟�Ud^���ڧ�G�h����F�)��fAr8㟫dNx$������7Gse˂����ntO?YP�N��Zyߚ�1O��ܤ�qf���	�&)껮}�Р���?�C:���ٵ�c��S}�a��U�6h_w�h(�����|ȹ\���$҉��'��8aXV���ؕ�RGŃ8?�봜��j����h����Ӗ�@ځ��$���E�P��V��+i�o���UYݎ�O �tH�>OJ�*���)�_o3 ����4�-Yj]�uMYԀ3��U�s�Q��k2�i�8;�߄h�՗��p��Pu"�{O?%|~�p7=���?�=�
�b���b1f��l5k�l�<�k�NIY������L�rM t8��t��m�2��J4�$6,�c|����t��
��.1*V���ܕ���D�>gs:F�m�-�6�l��V��}�����  ��/(�A��V�:ǖ�x���A�^�Q�GE���E�w��:HI��2��B|�#����p@�Z+���6	���JF�l0!l�I�B*
�D)��`��d���N�;��(�"|�5 ]|:����rª��� ұQ픡�����]6R���_��l��!���b^�=�\Q�/�6ȯL~cbU��V�*bM-�j��s�lq1�|u�s?���t]_� ��@�T?<CE��v�ݩ%Ӫ���.�!��;�/H�_��f�@D 0�?�u]��k��8O�l� �̈́�@��7� ��;r*[�0rR���^���Q�d&(�8;>*�iY���
΋���e�����?��+�"���ލ9Z%�oV
��,HRN(U�*e�rԃC�5�����+:�;?l_."�U�,�����f2ն���_����"�Cl��l)t}��0�t4`2���9Z��0��).�J�N�Гl�����HIp��晁��&M�j��k�]��^�e�cx�p�8RZFN�"|��{ńJH#P����QJ��{��Bzg��D�H���B�]ÀyX�ckJr:y1~Ğ�ī���%ɒ�5��d]f���� #�D#\�m�w�տ�v��Ze�Yn����KÙ��Q�L�^�n��W���h�R��<�!"c�7 @O����f�3��9��ٰ
6k� :ܽ�m�5/�a�E���c��X� �&�YpH�(�}�ȽND%x��B�F�v�k?�t�owqċD�0$�憰J�Աm�S�����;�����2uZHџ*jmp"��r:m���h�Œ&��3�*�\7��B�̣>nP9��0p,0x�t=Ȩ!!8�˖�c�:Poۑ"3��ऎ�J�Ge��Hܒ�:�=T��H?��5�h�����4��J��ƌ{�Y��3+��W�InLCN�w�w��Z��ە���D�zog����a�o���}���Ve*+����Bk��x_-Fd�T�|�yH�!W¾��i��@�V���KC�6�%��u�O���/�^���'x;GGu��!K#�y��ss!��Y���K\�h�|�7�T3����-�甌PjzZ���x�J�)�z��8k�o(�Tj��=�{�W&�f�n�G�#�7�Ρ�cRmuTЕ�sjv�jDA��;&��F�/���n*�e����;LYc���u��œ;뀍�
	�8)��U�C�����I�m�K�z����7�zj���X����5p�G
"��W��2�],�Ϭ=	�.�ݣR �až�J����Dv�F)$�Y���s�?>�Jiߵn���ͼ���
q�P��l�ݹ	d�����@�s�w4�/�"�n��D����4l�#lѸd�����eE =�ʷ���� t��S�)X�q�flk��-TL�I����ʁ�}�HU�_^#��Bs��w�<���{L}z5�G��:I�4N�5l��
�;ɍW=�z�ǐ�0Z�5G:A��b�U��領萷o%���'L�W݂�B�ڋ,!�3���s����Ʌ�yAl�B�r�,�P�z�-8]�(�ױH
q�s�O�L>e3gi[��U�h�.�e�����Y{��=N���7i
Iu�CY�b�&������!Rx(#�����&sG�.�/��^� '.PZ�T�W�t������2���;�@��x)��t���k-ו-�ˀobF�*Y���8���:�����4zV��Nt&2;>�ڕ�0�/Td�� `�
�9`~�zzfc�I0��D���y�JhP*�xrU�#��%'x��?��ٜ*�l@�)��Pe�`X�(z�ʸ��6y�I�����ֶ��8���ޓi�0z�O�N��q</d\3 �W4ub�!�$h�����5R�����7y	1���3'p����6m�[�'[�ɜ�A�o�FǑ�!����7�	s?s�ל�'V��'|N���f�O8.d5܀LU��Ox��~$�*޻�G���n~���<�-��5љh�|��ȩˮ 
ǋ�n�\�<]�
��9����vx�e��w̱��d�X� vd�!
ȵ�C\�U�3c����{��z)��q[�ܫ�����X��י�uw|�:���`�l^c3<؄��o4H�M{� �/R�tc��}��P��0s��U����]>^zCF��D��bD3�9Tw��cG�]�*�h�s��Z��a�#�N@5�Vۆ�q���^Cw����|����A���KΝ��:[���8����{�'�|.���<���8s����[���6�R��-�^�F��ہ��'F)�,�Ma��{��qs�B!�toz3�/M*�ߞI�Y��:WSjE�9<e�gOf� \���F�0�3�&Y�\��V8��I`)�+��(���=�k����a[��->Z�������`]٭�E�- ��Jի�H"�TB��ь15� EoLܧ|D� �^��X�C�6K��a�N������6-�bl������d�`�[=��LK���
A��w�
I6Ek�̯�p8��&�q�O�],�^+7�����C�>@=
�R�w`�\�A]B�	�!`�>���+���;i��W�ˤr���#B��R�gF`�a���1ni�q��*��6��\�(/ TX�:n=���g}3�.;��>u�VxNm_���l�@	Q>=�4���34�b���j��
_E���g`>S�z����b�(��P5��|ۭ�fM����`��6���S�l�a���0����^5B���:=	F7��������>٢��Z'�6O�Y�������Y�f�Ѝe����O��/3H�js�S7��������$�ﰰ\1�NدIg	��ty޴f�.5�o	����#_�a%��&�������x�챨P��~���|�gv1��+L���_!���w%#Z7P��7|,P������(F��}�t��	(-+&m��������͉��z�/1�`=�$���_�3{[mJ�)�.b�b�~��@��2��U�سQ�d��2srg�(�%�����j1❾��֥�r�R)f��)��wo�>�E�b�>���� �!�v�C{kv1ER��������=vå����������oa�Z��0J��5W��7��u�>��^M��|��IC Y^��䠰e��@�G������v��ܻʻgP|	8D]��d��/*�c=�n��9IzҞ�c���V����tȚ1�!�����das{v?��5��G\�T�t�5�I5qV�f�$�x�׌�(�Si����I�t6����t���;�ؖ?56�e�5]V��0+K�KxC�b��v����|lz��<��v��7�\�B�taTw٨�G�IAr�h�e{g��������J�s'�����Av/��U�R���c�
Ve���8s�bL Jtc%�sy��~�B�S1��X��lpT4�]�b[K؆���m¼^姫�ʚ+ar� �����\+K�eFH۸��yW�2��J� �����r�j9}�sgx$�?9���;/q��E�	B���%��u�(�ze���d�i3����XRQN��N:<�>A���������"���dB �)�f���������m�<CTm����%O�x�L0�c����26�_�F��}z �<y���\uU�r��#l܁���K)�T�>�Ճ�R�;?�-/@�$�U%����Ys9
���2��(�fl�L״��k;�a�Tg?�����*��.*��=k�%��-���~ܥ�w}�` �w��Ҙ�8���GB��?��Pm��D��蕟�M��S��e��/��@T�ۛ�77&�%e���βl�f(��>.�;��1���԰�QVuM)�h{�^<U��Y�e�N�f�V�.��f�����%�lDߺ����}t��+
Y��$�DM/�����F�c���g|�M����?)�gu7d�Z�+ �M�I��� ���P�E��S���x�2��I��@Rmx�/w�(Zg�s�������D��c��y�q{*(��>�N�X�_ӎD�偔��&�Y��,��䈩V&���N���2j��;+�,PH�[�pʹ���������Y��3r�ge�l���4Y:G��_ɗ�N݄����U��#��%,Ր�"˂�y>Fb�D��心���l���g�7�_F��u�of�[C���zi���ZK�\7ӭ�O�9w�<A%u���G��G*y��O�tK�}���T�<���*m3e;�dғ�d�U���z�1����2t��G�	Hݛ�(���$�˿������~x=wM�e8�8JZVue���m�1�av�Dv�����1�.%�=C�#�q�4t�P��WU���b �˥]w]"V�g��`a�lK@��;e�m��94�������b���������{�I��WV.�UR+�z�f���um���g3�-����X,C�w$�$	4��%�z7�IS9?��ۤ���M
�X�LځʉZI��0����H�GuU�j1��+3���a5G[&�Y$>"`q��d�Vj3�TK�UH@��~�Ȋ�'���~�)K��ωˬF�Uv�yʹ�ޘqܱ����gp��y��ߓ�>z��/�k�Ɛ�]@p6�I�+asO~<���1��P����[��{� �Y ?M ��#%�Ą�dq�=�`���<�g��[�����X{���c�1*H�"K.e�ҽW.�/�$FH��f��Z���7쁧��N�-��J2��Z�V:��0w ����]ߋ��R�TY���k-�@�bvJ����(Z��B!6�A��xw����9��t��\w�Ѽ�n{?4g+�ն�W�uX����,��`b	]'�l*.�e����
HN��	�<ߴ�s��[�c�$����L�^���*#!��̱�E�lA�3a�PO�,�����Ե�)�잼1��#e�9��<ٻ0���֠B֏]�=�� !�lK��`�ɕ?M3���Y�D�D-~��7pbw��-xUB��C,sb������ �\�6�����x1����v=&�p%�����&kQm�3�3sǨ�Z�
�.L ���84��|$R���F�÷��T���f�K�qJk��ZǴSf�n5t�T9&����-�F,�����t�.���H�"q�A�wu�F�)|���`ʸ�c��h��\�+��j�Q�aw����?F!�H�#7��x�L�=�a�4�V��3��*j`1�\E�����;?�����8�P{��Eu�)	�R��wD����T��D:�9�Q�2?i��f�M�<�3!�����X�Q%N��$�s�뀏IjM�� ��ah
�{S��k���=t�ߠ����ܦ��H�w�-a_<d�{�wm�Wt��ףt>�B7iF��S�����ALRMD@�!�-<Y\����Q���R�٥P��P�';�X.����� �ZBu�i��c�*^[�me��
����'g����1y��U<	��P�
��k����՛�����>8��E �j9`{�A�XU�������k���PF_�U ���T�I� ��; �<dl���C���+����eJ~��)��s�W���O��f�\"��r�	���R<�*�NQ���>P�.�5o}߮�QH��$�����0�C��Λ��:��m��d���F�b�*��Av*�p��Io�	�:�]"�:���v����5���������� �k���S�=ۏ!�z	�������4�Dwȣ�C+VIx��8��^��x�ZM��<sVg����a��߸N&OR�+��#	Ǘ-���P�3A8xҳ38�6o�GBMB�8#H�W��;f��Q@���e�T
[�O��t(���yR�'���(C1$"T�ni��l�t���s���Z�k�oC��_@״��	�&����Y7��z�n�v��v��0�D�-�r38����7%r�j�Jg���[ӺkcMj?q�v0�;��N�0E���H�L�^{٠�W�&#e�q���G�E���ʷ��Cr��ǈʤ��DK��X|jf�CF����|��xPY����_fL�>Ͽn�W�7��6���x1b��E<��@�z?��k��:��#�sM���6�4T��O.�1rԡ����
a2������,�E�J��2.�B��<x�o �4MZ�®$��`�/��Ty�;�c�����̢���rMn�p�x/忨��b�Z��_H� -yu@F%�O�NR4�5��I�^�
f��f�u%]|�u�b�\���u^�f��C)]tm�'��K��È�:-�G��a�}9�J^�h�I���1c�/�{���(�=�# O�3����]܀S1�(-	��=o�HQ��u�E	^x��)�e��I�8�<���x�-3��n�3��n�
T5l�NX*N�%������G��u����%}B��5#_�������31�i1�d���
v�}���9zu�n6wØy!�m#i�]����-�?J,���cx\��B�]m����$�������.Z�桅2A۽��P����{р*x(x�o� ���=?��%kD��[� ��bw,���(�_kʭ��m��U��T����ir�Zgh�)�[���s:m�%�%N�EO������_Q�7{���p����ZaZ�8i{��b6*bN�ji��r]+Yp�&<`��۱�3�%��>�4~�3�]ZtR�u�BM��%�Ue�^�!�D���ˎ>�XUU������E�U b`�в�
�n��A�����U�-��KEd��e�Ti�u~t�5N���z��R T���1��ޯl�kFy��&����J!y�:5p����'(!�c��CƔ�m�B=)yQ��#q7������)��Q�C^�M�����?��M��M�>�<hY�م9RP�N���2O+>�@��9��Y�rQQY��@Aw`Ո����d�[c$��FaB,�]�R�(���oef�c��[��6���5�8�_ι���e�w<R6ej:5�@=��T�~|�^�t���A�aoL���c�y�2GO<�����'�=��l��$��)V!���Yn��l+�ޑ�	0ˈ}�}:_�/��18Je�t�E k�֨N��債��W���Iq�����	�J��$��6-�AƸ�| ����T'�@9|d���$�HvC	xE�IK�׺k\�U�j?%g��q�Z��uL�O�&Iހ�Gga�"�����y�5�0WY��m�P��w��z�{�1fr���O�w�[L���k[���]�8�#j���I���+��g*H �Gpi�����ö-�u �.��m���0��5���$\q5��$�$<�А�:�2�/�x0J|�����":T���'e����s��W�ٹ�_�C\�x��`TŴ�F����;)X�Q����j�wH��������.Ljզ�h�B���-���>�(Gh_�Al=B���i5���j{\�k�'���T֌-�9lҼ<Υ�
�Z�v��gko�(n���Uf�?����4�1���߳lq�J"�ᄀ�C�j]��o.�(֌mQ/`��N\�j��g%(�9 ���Q�XV+�J�d�P�8�;�6�;��P���1?����H�N4+ugIԆV������۾���ʹ6�QPl�y��k��jx���
.sH_�g�.e0>#�w=q�w���j��e���ǳΤ�a6�%s��|��.nr�I�r��hm�u�X ;�2\(�����ZNe��d�!ͤ�)(ؕSd�xOC�L�' �|�OR�	� ݑ�����ۗ�'�J��q����}p8�q��П ���|w�5�D��0��m�����qkU�
t�5�������}8�^��|m!s������g�YZ���,�Ц�*����m~�΄�g��T��	�y1_�I�y	�Yǿ�P�5?� a>��("
�-kӈ�[ק�*���I�R��g�﫵���zQD�@s��
��z��|�m�����4Dgl�9Z�NV��\��bp�{#mZ�r���Q�x�w���k0h������Pt����󝖶C��yN�/��6w��l���Π�����;1d���%U�E��Մ�B����F�h@��V��0%���_���+����|�