��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D����gP�������������44��Pg��w�k�n�L�t�=�ʠ̲J�=�	�$tG�讧��p,��sC��Xu�_ S�	��mZK�qnu�*u"ǋ<�L*�2S���!��i�އh���
������)�=k��l��hx��I��} ���l��CaoK^G����F�HE���}�-���8���C��)�6v��q+���BɃ״��0�Ўl���Ax�`93Di�j�]��0x��uHo8ȁ�h�+���]�,L��uS��|�>5��9�8>�U̒ �|�o=���{�
'�[	��ԄgI.��Rs���Z�GݲB�_/h�_g�ˢGmYAa/E���,Ӥ`�΁b�d�@��+
��kz<ˤ(�w����0C݊��L87�C��������z��H�w��ڻJ�:>A��>I�B	�KW�-H��
 �ѶJ��;�\�16Ji�,�z}�:d�9E��_����Z���o-�[Ɯ��F$v�KG�%Z�:�oA4w�)[����:��z�X�o=B�e|�_2��ͰUSo����I#ظu��#x	oC}�v�%����KBU�2 p3 e�+�0ʝ��l�;$랉�A��t�h�?\�<��d"]���xuB�@3�{��e40/���GC��������ھΛ�HWR4��M�q��q��x�Gf�5�AW@{�-��LX�d��փ��Z�$�|�t��u�z(t�]7C�ua�Q�t��>l̘�9qaD���5:Ee��LsQ�����yEE����.]�����[�J	��o��)�	�V,�Ñ���+��3�Q��D�ʍJ^�"�q��F)���������Ү�'7�6�K<:�;��j�WKӉ���&�x�h��^J�4��j|mQ�p�A@����:�w����~�9�T�d_Z{؄� ��>h��g/gm>g����	q��Fu�D��,ͱ���h�R�����3ɣ�n�q߰U`MP}�ֶ�%� ���$�*l����%F����� R�J�a��t�ҢvF`A�Px �Ò�­���C�U���"�L�~�>�u��>����}��{A���������-��x��m����܆PFnh��Ȑ㟲�}=60���b\Q�s��]�*5��k����:u��W^�i�(�)�M���|U<��xC��'�(}�%��Udၤ���nǩ�����.1�N��y�/%I{W_��W�w��=%�u">Jn�g�^�������e(h�"C
Z:��^<oyF[#eB����_|���]Ll�����d.�4&��_<�`��4�d`��ğ҆�Y!�,��֠��1�y:&K5�ݴ6��Ofz�>:`��D? b�����Հ, ��1�;�G��
�'Ld��>3bT��/oӋ� �X�fu`�2Q����CM�n5��'��f/¤R�잽Ε�'���U�*;V�����D1��� �cfPqC,U�ܥ4(��8�'u��=ޏ�F�û3�:����C��ܲ���E˓�'���wp��X��O���y��,u��M�ڔ��&U�A���ͷ�6��p�
��V����/釣���ov6�K�)�e@k��G��);X�RƳ�)��8��dm_��i[�ŅQ��U�b���$H��l�R�]�J�\��ًFҠS����ݦ?دﶏ�,�{C�t�>�k�\��&�`t����~RA.�Ӳ ��/}D��W��NY�W���H]�]�7]%�|���>��U'��Ū�@^/��H�=e�-�,�� �|��6Mѷ���;U�G�����0v��.������^�v�N'����#}�Ǜaq6�HEc��i�A��g������ao���ޅN��-! �V �]��89�{��@�?!���KqK/�4X��qӦ�X7��n�5CӃχ���e��L�:Y}�y���(
�f8���Q5�?<r1��P�X[}�,"�44
�9y3�[Y�89�>����R�N��q�Һ���7�}i��$S����h:��^��\�9����ߚ��-�/�\j��Q��]
W����p�5}g��d�1�	{��W2^y���z�'�t�+�J|@|+`��mtqC嶁<u�$�
X���Ԯ���uW=;���EyF�C� �.��ƁI���,3�f����d�0 �T���-4����ʊ��:�(�$ �[i����ɸ��Qs^/��nBKtϨݺ��h�,Y�V�GSR�{?Y1�#�<nRץ�7�"�m�E��ዸmgJج1��]g�
��sm����E?|�����ꈛX����⻕A�2L�AC�Vh�u�n��P��o��C�Eu6c�}5��^^,dX$n/]7�u�XW/���]MDg�_����X	�U5�>T,��Q*E B��y9P�v[v�W>�F@�)��1{@��=ܑ������~�e���c�d��8�P~Ho1��aiivK���$���&�jc�I��%��v}�����N��;%����<�q��B������r��g��y�J��U5e�?I*���bD�ԫ6<o�s�lˮ��
�D�[O6J��Wt��	XK�����;7�^��d�'";dl�;0~h�<X�;U����sV|Ŕ���-@�1ʇH�m����|��X]��ۺ���\���b�^�G���VO�W+nN}�f��W{?�NQiCdX��2V��\���@\�Ȟ�aC�����LY��tԼ���n�F��p4� ��F�v�M��C&=��4��g\��)w����c��N�e{z㚆���KT�����sW�/�|6M!��c�Y�{�7L��J��5������5���vD;zڝ>��4H��9T�܌�(	���U�h#��K3��`j /���|L�0^��~�v����T�V�&�ql�w��c�UY�JpT4㨈h��'+k�?h-*M������X2?�g�Sb!���5̑���S����x��� X�T���=��f+&�,���� ~�[{�_N8��N���Ȝxr
��3�W^�Tt��7�Y�jH�MCd�g�ޡ�9��7����{�l�ی����Y�6ߏR����ҷ��&�WՄ�,k��I��H"͙�&�Z`F���7�i��V��cee�-%���)��u��q� J�Op��B�+ԥ /����dg
ȷ�p��IT�/]�n}���eRX]��@�%�8�����C_" �����x�A),ާ��'Ze{�ou,�M_v��)�o�֧�s�gDE�ޞ-=اJ�]��Y���1�,�
b�� ����:�����ż�H� ��] Q%RG?vG]���c����ܤ2vz.�BQF҂�jv���W|_K�n�뙱R��+S�-M6EVd[îH�ܨ7JSH�E^KC���cS�=�`�Vq���KZ_�p�B�8���O���V�ϹQ����Y��?R�Yڝ�##Hl�v��+��| e���Q��{�}5^�m����ջ3�d�b^E�\���zH��5�|ʤ(�,ޥ�*j6���Ҷ�F�v��Z�"9�r�}Bi� �Z�1*�;���3��\@{�O�ZW�Y�y�+�y���#`�L-r�o�8����/�����ؒ� ;��`��Pĸl_����P�jI���'q��K���W���z���i6�4�ԯ�1@�?����݄�L.�����{w��OaO%��_�	�$�-�����sX_e��]��:(�v^-h-�ne���BB⯛yO�>+09^ux���\k��B_�u���0�AyI��TP��L���0TM�����d���밊�0���!�\��	�5;8��vP5����ZT/�&��"�9ɍ����B�����^ԅ��z�/�_4�[�a��'�gK��a��)�uS����,c��{�B���6g࿦�O���b��&y�V�V�K��z�gw�\���.����P'�n@��n��M��9y�M��!ym���cѱ,��LCj[�P%۱�J��
U:IQ��Ry���0�B�L�xegL�*a����%�:S�G���pF�J)���sQBɌ�G�1�T1�[4�tʀ+�*�t��RR�s���{F q��"��|�a	�[��@�&A`��]'8P�qv��Bjh�{Ő�/P�T��ь�2M���ә��;�fB �ZIu��x�:K��B0� �U�%��l)�vj��y;$`l���[��`>K+LZ�쿫)��P}�4	~��SЯt<������>�PE�������l�VѸ$c>M�JY���i�\����E �";< ����"�����#{���������W��AL_>���	o�.oq������?^��6���#��~�,P�cڴv���<� ��1�P'�/y3=7�|`b�03�Q����EUV��g�E��cW�ULù�r����x*ux�Q&��� Y���4 ;F�R#;*�U�XՃ �2��ϒ"qnP��;ڲ���s�O��ůP�#U��@a� "�M7h��vyr��L7:��8�In�U
.�5��1=;B���.�my�~��8�[jy}�k����=�y�'}M��E�P6A�g=
=�cQ���j�{�ļc��p4��9[%�^3$���4[��lUu
��\��8�M���׺>�o����jU����9(�5qńB9l��Lަ�.}���@t{t�w0��v�5�O6v-[n�l��}��夵v��F����\�a���r�j6/���`�^�^��kV��x�$ ���R�/h'�	���h�t�c)P��V�s'\.���J�汽s�2���/z>S���۽l�,�͕j�H���QȒl��e'
�VJڊ斊7-$m}�)�Kٗk�0{�����i��^D�\ ���|4��v�i\�˧	v��0Tb�ޟ�u���N�6B��P�M���Ɨ�/�W�XiW�T�!�G�����g'7�<j�{��4�C�b�⊝��@2����i�*''p�2��s�g�g�\2;:���?c�ԑ�V��NI��u�; �&�r��a��St���-����(\����c�K�úz�����5���o²V9iJ���櫉�Er��.MZ�De�6��h�f��<^����U��"����k}�TY�ig��dD	R�@���A�GHuX�tx�����7,�ab�s7�!0��҈_潦5G=�bk��ҿ^*�z5���,cs匬��f�Q:�+�g�e,��(�;}��Go]���&R�П(��!�\AzgAN�ͣŕC��W���Q�Cӟ�K��}h�J��������ڨ�0��ʋׯ��%��/%���w�=�,���?��dX"4��_��������?�?�do�E�ۥr�OKe���9�O\7?��?�A�tqְj�ʜ��Y�$d�r��ygͦ��R�E��[d��+�7)׸���SCk��7�4�0�<���� �`: �nhyG3����~~�׫�>kd�X�B��l��
qT 7�H
���ؑ�OfEj�~�������������s���0)knU���F2�<`�Y�,n��q_G�J�ڤz������A���W�Á���k��x��abt�+����;Nڏ[�:�&��t�O�K��Ҵ=�e�|H�J�Y��Ň�'��ަlQ��~m6��z�Tr
�ɱ-��B���z�&���x�J�Ӭ�`�/�E'���3�J4-����#0�c�h°�bZ
�m�����QuE�A��%o��n�8���ٝ)Si-�r`!m	�����?�jZ��T
V�*��k����ó��n �8 �> � ��l�q!���2jl����?D��؞�,!)ߨQu�dP6$X�RJ�Up��0�(k��Y�^Γ)�U�۳����(^˺��e�wg_fA_��F�
vܙ8�00!L�Y%ci\�"7���@�'� ����'���:M��ux�h�����T'vP�`��8���-рO�8����y�>O����r'�9�\��5���\�z�ٮ]^�q�b�OB\�ėҤ�]��;����j��r?�p܍��)��[����r*o���ܕ'�#j�[�M���rnE ��AG\=G��@���$�`���SHV;qtW�sTp�9�/���)>(&��n<����p(�X㲞�Q��b���dmHM8��I⨔�׊9
n]I���Ae�9�v�3�ƚ���VJ~�v[/"���lq��t2Qa]�χ�� �U� ѳ��Ҥ��=�������T3,����}И�uB�z�hD���+eIq]�0lX_�5'�q�]U�f6#k�|��U���剃�SGN`�ڲB1뱽�+�I��z�1�xJ��WH�<�γ������ �F�'PqG?����bzڊ1�Z(��O[l
Jyq��`��:�[#�0&�|�PM1�)����;~�|Mغ��V�RO
:\F�^��*�(a���3���w�J<O�C��)O����"��F����ls)�3^��X�*��YL�,���F�9�o��?�]t�� �if*��eF��X�X!���쮓v���Q�Z�E���-�oKt��K�`|u��mb ���g�gi����=��gͮE��i��>ZO���&=���׸��٠B2�����'L|G���WʍƨT̌m?7ܬz�V2oֈ&�sw�'�A��_���0��q�U��w�Y���\���2R�Wxk E
���ȯJ=no�p�5"���M�P/�W�\UJ�=o��:�1u��	�=ց�7ze�1�[�s5�4��r�Ld����*�R(fC�E ��U�c��n&�jm�Vr��I�]o��R�nω�=R�L�#	��46;�Ni�k�Y�c�G�3U�LH��b�G	����t�,5�	Tb8�����cuߜ��1%G�J�`?�y�ٴ~��.˪+#��%�T�Q�N�̬oy�|��K��p��*\�0���� Ͳ���SsP�c(@�H��s��ID)�d
w��}5���iUQ���H�K�,���F��fA"+%�e�%7zT��}!�1?�4�z(:�LT�v��R&��~���8�S)՝�	���������9v�_~��ݎ.e�8�m�]�0����q��]=�(��0�|j4V]3�*B!�f̒^��!�^ZJhȗ�7iU�� �A6�ߊ���k�a��^�_d~�3��J+ "$T��HP��ۯ�kb�e���/����H�8#Iu��rf�'BM"���M��0cC�c����އ~�[$3�r��&��n���);	IvN�ټK����<\MAd�[�e��Euf��r>!3�_wUI,~Y1�)x8+4���X��ݠJ�|u@5�r�-Vs�At�_(2�^���9��_��Ǖ$ t,u���(�O&�C\���p���h�"���SGGMyjf����K������b���rT�x<� �L�4k]ݣ�h��櫁��"z԰`�Z��cT�Y~ڋ��ś|yG_"�P���/��vJ��W��Z@';7����+�����"�>���;^��,*������-vnXv���"�,�P�)k��w�r�^���j-T����\جG�횔�� ےKvz�(i���X��:wh#v�����:�m0e�mo_;�����KS⬃�4�`D�O��)I�l(\r��$�2T�AE���`��ޣ�������f�H����#�s��ɬz"]���,��1o�� ��j��_<�ft@f��z`�-{9�d���iܣ���y�����H������9웆��}�݂,�<�Zʢy��ue1�[�B޺��b+��t�q G�D���e�W�j��i-c��7�bp�HKM��P�O��m����M�����ԁ�`����'���MXnd��
�������M> ؜��5����^pA.��pY��$ev�����/�Щ�E��f^Gg�]�۞���+�d���N�/n
Ĵ4��S>��w3wAK�a�&�(����-�+Kc��׌[e�����rQ|f1X9����~��Ÿ�;-��ƒ��A��C��[�D��GP�����`�J�]����H�9�;�=Z�2��	,��=��؁A�Y�]�.�뮸���f�c��g:�Ō'h��8��4CM�#�#!1� h��!k��>�Iro!�7H�/�c*}W�uyײ��g�p�mH,U(��X��<��L�ܳs@�w����۝�f:��ƶv�K��z�����;`���4.6�����kZ?B��_<���̘�nU��e�^��/����K��Z��b�4��{Cu5ޚ��XL�����H��aۚ�4�p"��qX��EMFCf��fD��i4	0�`2��������d	A�P����^X*�xq^�����a5iĸ�#�S�hT�b�`w��?��Hv	׏��?�^��Y7~�����[���ƴZo]����7�do�-A�߳=.�3n��ᜅ��{��� ��:��6�Q����q��������GN�UWw�i����sM�:Ľ�Bj�s`#���c܍!K0p��q��e�6m6WQ|�$[���Hڨ�+$�ϖ����Մ^:�y��	I0����M����t>�eV����JΊ����ڜ�"9X,	#:��]M��\C���U�8��-�=��u8X�|�S��	Iڸ#⯦^N��