library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

entity console_glyphrom is
    port (
        clk : in std_logic;
        address : in std_logic_vector(7+4 downto 0);
        din : in std_logic_vector(7 downto 0);
        dout : out std_logic_vector(7 downto 0);
        we : in std_logic
    );
end;

architecture RTL of console_glyphrom is
    type RAM_TYPE is array (natural range <>) of std_logic_vector(7 downto 0);
    subtype BRAM_TYPE is RAM_TYPE(0 to 2 ** (8+4) - 1);

    signal BRAM : BRAM_TYPE := (
        x"00", x"00", x"7E", x"42", x"42", x"42", x"42", x"42", x"42", x"42", x"42", x"7E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"7C", x"82", x"AA", x"82", x"82", x"BA", x"92", x"82", x"82", x"7C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"7C", x"FE", x"D6", x"FE", x"FE", x"C6", x"EE", x"FE", x"FE", x"7C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"6C", x"FE", x"FE", x"FE", x"FE", x"7C", x"38", x"10", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"10", x"38", x"7C", x"FE", x"7C", x"38", x"10", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"10", x"38", x"38", x"10", x"54", x"FE", x"FE", x"54", x"10", x"38", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"10", x"10", x"38", x"7C", x"FE", x"FE", x"7C", x"10", x"10", x"38", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"3C", x"3C", x"18", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"E7", x"C3", x"C3", x"E7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"24", x"24", x"18", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"E7", x"DB", x"DB", x"E7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", --
        x"00", x"00", x"1E", x"06", x"0A", x"12", x"38", x"44", x"44", x"44", x"44", x"38", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"38", x"44", x"44", x"44", x"44", x"38", x"10", x"7C", x"10", x"10", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"3E", x"22", x"3E", x"20", x"20", x"20", x"20", x"20", x"20", x"C0", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"7E", x"42", x"7E", x"42", x"42", x"42", x"42", x"42", x"42", x"44", x"80", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"10", x"92", x"54", x"38", x"EE", x"38", x"54", x"92", x"10", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"C0", x"F0", x"FC", x"FF", x"FC", x"F0", x"C0", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"03", x"0F", x"3F", x"FF", x"3F", x"0F", x"03", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"10", x"38", x"54", x"10", x"10", x"10", x"10", x"54", x"38", x"10", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"24", x"24", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"7E", x"92", x"92", x"92", x"92", x"72", x"12", x"12", x"12", x"12", x"00", x"00", x"00", x"00", --
        x"00", x"38", x"44", x"40", x"30", x"48", x"44", x"44", x"24", x"18", x"04", x"44", x"38", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"7E", x"7E", x"7E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"10", x"38", x"54", x"10", x"10", x"10", x"54", x"38", x"10", x"7C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"10", x"38", x"54", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"54", x"38", x"10", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"08", x"04", x"FE", x"04", x"08", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"20", x"40", x"FE", x"40", x"20", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"40", x"40", x"40", x"40", x"40", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"24", x"42", x"FF", x"42", x"24", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"10", x"10", x"38", x"38", x"7C", x"7C", x"FE", x"FE", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"FE", x"FE", x"7C", x"7C", x"38", x"38", x"10", x"10", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"00", x"10", x"10", x"00", x"00", x"00", x"00", --
        x"00", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"24", x"24", x"24", x"7E", x"24", x"24", x"7E", x"24", x"24", x"24", x"00", x"00", x"00", x"00", --
        x"00", x"10", x"10", x"7C", x"92", x"90", x"90", x"7C", x"12", x"12", x"92", x"7C", x"10", x"10", x"00", x"00", --
        x"00", x"00", x"64", x"94", x"68", x"08", x"10", x"10", x"20", x"2C", x"52", x"4C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"18", x"24", x"24", x"18", x"30", x"4A", x"44", x"44", x"44", x"3A", x"00", x"00", x"00", x"00", --
        x"00", x"10", x"10", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"08", x"10", x"20", x"20", x"20", x"20", x"20", x"20", x"10", x"08", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"20", x"10", x"08", x"08", x"08", x"08", x"08", x"08", x"10", x"20", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"24", x"18", x"7E", x"18", x"24", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"10", x"10", x"7C", x"10", x"10", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"10", x"20", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"10", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"04", x"04", x"08", x"08", x"10", x"10", x"20", x"20", x"40", x"40", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"3C", x"42", x"42", x"46", x"4A", x"52", x"62", x"42", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"08", x"18", x"28", x"08", x"08", x"08", x"08", x"08", x"08", x"3E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"3C", x"42", x"42", x"02", x"04", x"08", x"10", x"20", x"40", x"7E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"3C", x"42", x"42", x"02", x"1C", x"02", x"02", x"42", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"02", x"06", x"0A", x"12", x"22", x"42", x"7E", x"02", x"02", x"02", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"7E", x"40", x"40", x"40", x"7C", x"02", x"02", x"02", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"1C", x"20", x"40", x"40", x"7C", x"42", x"42", x"42", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"7E", x"02", x"02", x"04", x"04", x"08", x"08", x"10", x"10", x"10", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"3C", x"42", x"42", x"42", x"3C", x"42", x"42", x"42", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"3C", x"42", x"42", x"42", x"42", x"3E", x"02", x"02", x"04", x"38", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"10", x"10", x"00", x"00", x"00", x"10", x"10", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"10", x"10", x"00", x"00", x"00", x"10", x"10", x"20", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"04", x"08", x"10", x"20", x"40", x"20", x"10", x"08", x"04", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"7E", x"00", x"00", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"40", x"20", x"10", x"08", x"04", x"08", x"10", x"20", x"40", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"3C", x"42", x"42", x"42", x"04", x"08", x"08", x"00", x"08", x"08", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"7C", x"82", x"9E", x"A2", x"A2", x"A2", x"A6", x"9A", x"80", x"7E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"3C", x"42", x"42", x"42", x"42", x"7E", x"42", x"42", x"42", x"42", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"7C", x"42", x"42", x"42", x"7C", x"42", x"42", x"42", x"42", x"7C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"3C", x"42", x"42", x"40", x"40", x"40", x"40", x"42", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"78", x"44", x"42", x"42", x"42", x"42", x"42", x"42", x"44", x"78", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"7E", x"40", x"40", x"40", x"78", x"40", x"40", x"40", x"40", x"7E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"7E", x"40", x"40", x"40", x"78", x"40", x"40", x"40", x"40", x"40", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"3C", x"42", x"42", x"40", x"40", x"4E", x"42", x"42", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"42", x"42", x"42", x"42", x"7E", x"42", x"42", x"42", x"42", x"42", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"38", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"38", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"0E", x"04", x"04", x"04", x"04", x"04", x"04", x"44", x"44", x"38", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"42", x"44", x"48", x"50", x"60", x"60", x"50", x"48", x"44", x"42", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"7E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"82", x"C6", x"AA", x"92", x"92", x"82", x"82", x"82", x"82", x"82", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"42", x"42", x"42", x"62", x"52", x"4A", x"46", x"42", x"42", x"42", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"3C", x"42", x"42", x"42", x"42", x"42", x"42", x"42", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"7C", x"42", x"42", x"42", x"42", x"7C", x"40", x"40", x"40", x"40", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"3C", x"42", x"42", x"42", x"42", x"42", x"42", x"42", x"4A", x"3C", x"02", x"00", x"00", x"00", --
        x"00", x"00", x"7C", x"42", x"42", x"42", x"42", x"7C", x"50", x"48", x"44", x"42", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"3C", x"42", x"40", x"40", x"3C", x"02", x"02", x"42", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"FE", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"42", x"42", x"42", x"42", x"42", x"42", x"42", x"42", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"42", x"42", x"42", x"42", x"42", x"24", x"24", x"24", x"18", x"18", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"82", x"82", x"82", x"82", x"82", x"92", x"92", x"AA", x"C6", x"82", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"42", x"42", x"24", x"24", x"18", x"18", x"24", x"24", x"42", x"42", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"82", x"82", x"44", x"44", x"28", x"10", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"7E", x"02", x"02", x"04", x"08", x"10", x"20", x"40", x"40", x"7E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"38", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"38", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"40", x"40", x"20", x"20", x"10", x"10", x"08", x"08", x"04", x"04", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"38", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"38", x"00", x"00", x"00", x"00", --
        x"00", x"10", x"28", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"00", x"00", --
        x"10", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"3C", x"02", x"3E", x"42", x"42", x"42", x"3E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"40", x"40", x"40", x"7C", x"42", x"42", x"42", x"42", x"42", x"7C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"3C", x"42", x"40", x"40", x"40", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"02", x"02", x"02", x"3E", x"42", x"42", x"42", x"42", x"42", x"3E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"3C", x"42", x"42", x"7E", x"40", x"40", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"0E", x"10", x"10", x"7C", x"10", x"10", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"3E", x"42", x"42", x"42", x"42", x"42", x"3E", x"02", x"02", x"3C", x"00", --
        x"00", x"00", x"40", x"40", x"40", x"7C", x"42", x"42", x"42", x"42", x"42", x"42", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"10", x"10", x"00", x"30", x"10", x"10", x"10", x"10", x"10", x"38", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"04", x"04", x"00", x"0C", x"04", x"04", x"04", x"04", x"04", x"04", x"44", x"44", x"38", x"00", --
        x"00", x"00", x"40", x"40", x"40", x"42", x"44", x"48", x"70", x"48", x"44", x"42", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"30", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"38", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"FC", x"92", x"92", x"92", x"92", x"92", x"92", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"7C", x"42", x"42", x"42", x"42", x"42", x"42", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"3C", x"42", x"42", x"42", x"42", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"7C", x"42", x"42", x"42", x"42", x"42", x"7C", x"40", x"40", x"40", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"3E", x"42", x"42", x"42", x"42", x"42", x"3E", x"02", x"02", x"02", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"5E", x"60", x"40", x"40", x"40", x"40", x"40", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"3E", x"40", x"40", x"3C", x"02", x"02", x"7C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"10", x"10", x"10", x"7C", x"10", x"10", x"10", x"10", x"10", x"0E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"42", x"42", x"42", x"42", x"42", x"42", x"3E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"42", x"42", x"42", x"24", x"24", x"18", x"18", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"82", x"82", x"92", x"92", x"92", x"92", x"7C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"42", x"42", x"24", x"18", x"24", x"42", x"42", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"42", x"42", x"42", x"42", x"42", x"42", x"3E", x"02", x"02", x"3C", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"7E", x"04", x"08", x"10", x"20", x"40", x"7E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"0C", x"10", x"10", x"10", x"20", x"10", x"10", x"10", x"10", x"0C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"30", x"08", x"08", x"08", x"04", x"08", x"08", x"08", x"08", x"30", x"00", x"00", x"00", x"00", --
        x"00", x"62", x"92", x"8C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"10", x"28", x"44", x"82", x"82", x"82", x"82", x"FE", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"3C", x"42", x"42", x"40", x"40", x"40", x"40", x"42", x"42", x"3C", x"10", x"10", x"20", x"00", --
        x"00", x"00", x"24", x"24", x"00", x"42", x"42", x"42", x"42", x"42", x"42", x"3E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"08", x"10", x"00", x"3C", x"42", x"42", x"7E", x"40", x"40", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"18", x"24", x"00", x"3C", x"02", x"3E", x"42", x"42", x"42", x"3E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"24", x"24", x"00", x"3C", x"02", x"3E", x"42", x"42", x"42", x"3E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"10", x"08", x"00", x"3C", x"02", x"3E", x"42", x"42", x"42", x"3E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"18", x"24", x"18", x"3C", x"02", x"3E", x"42", x"42", x"42", x"3E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"3C", x"42", x"40", x"40", x"40", x"42", x"3C", x"10", x"10", x"20", x"00", --
        x"00", x"00", x"18", x"24", x"00", x"3C", x"42", x"42", x"7E", x"40", x"40", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"24", x"24", x"00", x"3C", x"42", x"42", x"7E", x"40", x"40", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"10", x"08", x"00", x"3C", x"42", x"42", x"7E", x"40", x"40", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"48", x"48", x"00", x"30", x"10", x"10", x"10", x"10", x"10", x"38", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"30", x"48", x"00", x"30", x"10", x"10", x"10", x"10", x"10", x"38", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"20", x"10", x"00", x"30", x"10", x"10", x"10", x"10", x"10", x"38", x"00", x"00", x"00", x"00", --
        x"24", x"24", x"00", x"3C", x"42", x"42", x"42", x"7E", x"42", x"42", x"42", x"42", x"00", x"00", x"00", x"00", --
        x"18", x"24", x"18", x"3C", x"42", x"42", x"42", x"7E", x"42", x"42", x"42", x"42", x"00", x"00", x"00", x"00", --
        x"08", x"10", x"00", x"7E", x"40", x"40", x"40", x"78", x"40", x"40", x"40", x"7E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"6C", x"12", x"72", x"9E", x"90", x"90", x"6C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"7E", x"90", x"90", x"90", x"FC", x"90", x"90", x"90", x"90", x"9E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"18", x"24", x"00", x"3C", x"42", x"42", x"42", x"42", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"24", x"24", x"00", x"3C", x"42", x"42", x"42", x"42", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"10", x"08", x"00", x"3C", x"42", x"42", x"42", x"42", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"18", x"24", x"00", x"42", x"42", x"42", x"42", x"42", x"42", x"3E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"10", x"08", x"00", x"42", x"42", x"42", x"42", x"42", x"42", x"3E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"24", x"24", x"00", x"42", x"42", x"42", x"42", x"42", x"42", x"3E", x"02", x"02", x"3C", x"00", --
        x"24", x"24", x"00", x"3C", x"42", x"42", x"42", x"42", x"42", x"42", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"24", x"24", x"00", x"42", x"42", x"42", x"42", x"42", x"42", x"42", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"10", x"10", x"7C", x"92", x"90", x"90", x"90", x"92", x"7C", x"10", x"10", x"00", x"00", --
        x"00", x"00", x"18", x"24", x"20", x"20", x"78", x"20", x"20", x"20", x"22", x"7E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"82", x"82", x"44", x"28", x"10", x"7C", x"10", x"7C", x"10", x"10", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"F0", x"88", x"88", x"88", x"F4", x"84", x"8E", x"84", x"84", x"82", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"0C", x"12", x"10", x"10", x"7C", x"10", x"10", x"10", x"10", x"10", x"10", x"90", x"60", x"00", --
        x"00", x"00", x"08", x"10", x"00", x"3C", x"02", x"3E", x"42", x"42", x"42", x"3E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"08", x"10", x"00", x"30", x"10", x"10", x"10", x"10", x"10", x"38", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"08", x"10", x"00", x"3C", x"42", x"42", x"42", x"42", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"08", x"10", x"00", x"42", x"42", x"42", x"42", x"42", x"42", x"3E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"32", x"4C", x"00", x"7C", x"42", x"42", x"42", x"42", x"42", x"42", x"00", x"00", x"00", x"00", --
        x"32", x"4C", x"00", x"42", x"42", x"62", x"52", x"4A", x"46", x"42", x"42", x"42", x"00", x"00", x"00", x"00", --
        x"00", x"38", x"04", x"3C", x"44", x"3C", x"00", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"38", x"44", x"44", x"44", x"38", x"00", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"10", x"10", x"00", x"10", x"10", x"20", x"42", x"42", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"7E", x"40", x"40", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"7E", x"02", x"02", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"20", x"60", x"20", x"22", x"24", x"08", x"10", x"20", x"4C", x"92", x"04", x"08", x"1E", x"00", x"00", --
        x"00", x"20", x"60", x"20", x"22", x"24", x"08", x"10", x"22", x"46", x"8A", x"1E", x"02", x"02", x"00", x"00", --
        x"00", x"00", x"10", x"10", x"00", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"12", x"24", x"48", x"90", x"48", x"24", x"12", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"90", x"48", x"24", x"12", x"24", x"48", x"90", x"00", x"00", x"00", x"00", --
        x"88", x"22", x"88", x"22", x"88", x"22", x"88", x"22", x"88", x"22", x"88", x"22", x"88", x"22", x"88", x"22", --
        x"AA", x"55", x"AA", x"55", x"AA", x"55", x"AA", x"55", x"AA", x"55", x"AA", x"55", x"AA", x"55", x"AA", x"55", --
        x"EE", x"BB", x"EE", x"BB", x"EE", x"BB", x"EE", x"BB", x"EE", x"BB", x"EE", x"BB", x"EE", x"BB", x"EE", x"BB", --
        x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", --
        x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"F0", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", --
        x"10", x"10", x"10", x"10", x"10", x"10", x"F0", x"10", x"F0", x"10", x"10", x"10", x"10", x"10", x"10", x"10", --
        x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"E8", x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"28", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"28", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"10", x"F0", x"10", x"10", x"10", x"10", x"10", x"10", x"10", --
        x"28", x"28", x"28", x"28", x"28", x"28", x"E8", x"08", x"E8", x"28", x"28", x"28", x"28", x"28", x"28", x"28", --
        x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"28", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"08", x"E8", x"28", x"28", x"28", x"28", x"28", x"28", x"28", --
        x"28", x"28", x"28", x"28", x"28", x"28", x"E8", x"08", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"10", x"10", x"10", x"10", x"10", x"10", x"F0", x"10", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", --
        x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", --
        x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"1F", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"FF", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", --
        x"10", x"10", x"10", x"10", x"10", x"10", x"1F", x"10", x"1F", x"10", x"10", x"10", x"10", x"10", x"10", x"10", --
        x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"2F", x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"28", --
        x"28", x"28", x"28", x"28", x"28", x"28", x"2F", x"20", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"20", x"2F", x"28", x"28", x"28", x"28", x"28", x"28", x"28", --
        x"28", x"28", x"28", x"28", x"28", x"28", x"EF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"EF", x"28", x"28", x"28", x"28", x"28", x"28", x"28", --
        x"28", x"28", x"28", x"28", x"28", x"28", x"2F", x"20", x"2F", x"28", x"28", x"28", x"28", x"28", x"28", x"28", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"28", x"28", x"28", x"28", x"28", x"28", x"EF", x"00", x"EF", x"28", x"28", x"28", x"28", x"28", x"28", x"28", --
        x"10", x"10", x"10", x"10", x"10", x"10", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"10", x"10", x"10", x"10", x"10", x"10", x"10", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"28", --
        x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"10", x"10", x"10", x"10", x"10", x"10", x"1F", x"10", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"10", x"1F", x"10", x"10", x"10", x"10", x"10", x"10", x"10", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"28", --
        x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"FF", x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"28", --
        x"10", x"10", x"10", x"10", x"10", x"10", x"FF", x"10", x"FF", x"10", x"10", x"10", x"10", x"10", x"10", x"10", --
        x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", --
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", --
        x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", --
        x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", --
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"3A", x"46", x"44", x"44", x"44", x"46", x"3A", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"38", x"44", x"44", x"48", x"7C", x"42", x"42", x"42", x"42", x"7C", x"40", x"40", x"40", x"00", --
        x"00", x"00", x"7E", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"7E", x"42", x"42", x"42", x"42", x"42", x"42", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"7E", x"40", x"20", x"10", x"08", x"08", x"10", x"20", x"40", x"7E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"3E", x"44", x"44", x"44", x"44", x"44", x"38", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"42", x"42", x"42", x"42", x"42", x"46", x"7A", x"40", x"40", x"40", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"FE", x"10", x"10", x"10", x"10", x"10", x"0C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"10", x"7C", x"92", x"92", x"92", x"92", x"92", x"92", x"7C", x"10", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"3C", x"42", x"42", x"42", x"5A", x"42", x"42", x"42", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"3C", x"42", x"42", x"42", x"42", x"42", x"42", x"24", x"24", x"66", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"3E", x"10", x"08", x"3C", x"42", x"42", x"42", x"42", x"42", x"3C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"7C", x"92", x"92", x"92", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"02", x"04", x"7C", x"8A", x"92", x"92", x"A2", x"7C", x"40", x"80", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"1E", x"20", x"40", x"7E", x"40", x"20", x"1E", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"3C", x"42", x"42", x"42", x"42", x"42", x"42", x"42", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"7E", x"00", x"00", x"7E", x"00", x"00", x"7E", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"10", x"10", x"7C", x"10", x"10", x"00", x"7C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"20", x"10", x"08", x"04", x"08", x"10", x"20", x"00", x"7C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"04", x"08", x"10", x"20", x"10", x"08", x"04", x"00", x"3E", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"0C", x"12", x"12", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", --
        x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"90", x"90", x"60", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"10", x"10", x"00", x"7C", x"00", x"10", x"10", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"32", x"4C", x"00", x"32", x"4C", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"18", x"24", x"24", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"06", x"04", x"04", x"04", x"04", x"44", x"44", x"44", x"24", x"14", x"0C", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"38", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"18", x"24", x"04", x"08", x"10", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"3C", x"3C", x"3C", x"3C", x"3C", x"3C", x"00", x"00", x"00", x"00", x"00", --
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00" --        
    );
    signal ad_w, ad_r : integer range 0 to 2 ** 8 - 1;

begin

    ad_w <= conv_integer(address);

    process (clk) begin
        if (clk'event and clk = '1') then
            if (we = '1') then
                BRAM(ad_w) <= din;
            end if;
            ad_r <= ad_w;
        end if;
    end process;

    dout <= BRAM(ad_r);

end;