��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�Tں~�ImW�.�^�ᆹ��������]��%�wx����xeՍ�ϡ�&JLc7e��~�'[�b(�Z��M%기_��H�K%_N�kV�.���a�����F����B�u�E�[�D��*{2<(ڡ�Ki;�e��W�*�]�?eey�J�Agm��^��F�}��!kw���Ȥ�|m�B�9�Y{F�G#��=���]�q�x�>�dO��&���U �XF������[�K���b�h�s�����61�QSt���E�������Ec�,��t6�p4�%�&sg(s=��R*�iGHdIWr6���^�9�v})�X���m����ie�.7�~n�|p�=&��H�%��5"���*��K.Fhg�X�b�F�*6r>��Y�.���V����cH.<��#�I�;�'δ���}Z�gs�q����Hm��Dg�+����H��_�#QӴ!ͻ����w��l���zl|䎾m�Ի�G ����{���o�<,�[�f�1�j��/��L��X����0o[Ln�>O�l��~��E�V��(A�5��%1���u�n4c@a�!���5z�DE�{���8�Ƅ�xh����{'�pȘa$��B�i>g@������$��fud�6�7���i��mθY�N�y��G�tm7,���	�����f;W��E�����n0q]f�/v�oK���}3��Y�y6���p�M���a�z�j�xG��Kw��j ���$�'���_�]��z[qӡ�
�_�-.A|B�h�֫�3h!��
Z�:'��ډ�Cg����z_1ch�@���O&��ɤ�Y�����7ktL�������v=�M�'�/������,ŢL9�`8��EWo�)m�Y�R���@T�����-.O^Q!u���oR�6��n�Z	<�~%��o���?kD�ٺmTQ��Z���:�=:���^�L6p�~�4��9rK^J�P�^a�I�R��HgP�<��l��U��H&�'��9�Ĩ�F�|���OиsgβVf�$���UKIC�����U��[$��{���w��i��[�PA���b<��Z����߿VmU�~�d����'���P�_�L���m#j��"��X[+/NZRbtv�;�O�ǚ�,,�
�`=&���X�_5�5��u}���El���I���N%�A	я&7�R�z���E٢�uY	�0sI���Y�n��u#�m��3�p2Q��q�?\D�?l��6����U���nN����_��A�:(����1�'Q����9c�&�ג��@�w>�fH�B��]��}j�D`,�C��P9�U/|;%��)��}xeU��6DΠA��φ���z�ڿ��E���'�ӣ�Z���Wa�Y;�2�J�@��?���>�d��H�O���jvh��o�b����|Pl�����J���F��d�j���Y��g�U`/�1�C�U~�F�K�M%�(Z�I�L8��z;+�,P�/��0zX�3���C��֜�V�����;gﾦd�F�T�9u����f��R���<���(�V#�y��?�']��æT�Αx��윬�/3��r�<ۻ���[��֛%����Kvy[��#LA�	��<F�>M��rAb�!ڀ�u%߉�q"�[R�:����I8,5�!x