��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��5�����E�V��B�45�H]"M}�"=U<D���فlQ��Mn���d�Y�Σ14��V����y)��>]΄�F�Q0.���=�SF;��Ǉu���'n�y8���r�b-�I��7"/����/q�{Y(����P�bA�b�<�E?U��F:��f����Ki��;��i<��]|S�5���+����l/�vD������d���=F����v6L��o�S�����AgA��W��f�������e����+�ٯއ�%F7�8|K����^�0��o��A{��O�_���`�Qy��Us˩���i�6���?
�<�i"sě%5��Y7e�i�Y��H_��X�B������a��B|��u�cT2.�){�ê9n/ڭ�ZﾹH�Y�����C-Y(&Q�/
�
��}_`v�J��J��!�	r��9�Ea��	kQH�G=xXz��%��DP�!����<$�P����� ��J��bxhS��nr|�B����_�ʰ$f1I�D}��*�g��[n��U��S33؀�U�C� ����UȬ�����=�	)�`�*RI�0i��h�� �}`J7�%S���a:��+��C}e��w�v�������l1�ڧ�+��w�/�}����k���=�
�?���ø�^Ht�O��sf�XcI.��2�]���j��k\#x�<�hʺ*g�9�����@�
	��'"���1qA���m�L�U�8KG�DzC�4l,+�Qa]�B��u�{�i`���<1������������K����������Mq�� q'#�ʡ͏V��Sۺ�m���7��֪�C޹ ��Z��#1�t!K๝�I,�>5�qV��#L@��I�:.,{����*�	��L%k�̿����@����q�lx��-<��K�����c�)@j��")���������b�	�Ўg�=�*0����2}�0��R�-�?��eŽ��!���T��e�=�B�+�Z�Ÿ���S�O�ԓ�4ĉ�5��x0\{��|��F�΅7�pp*��![}�~��uZS�?i���~������|��8��@6xd�����eh�/��� �"
r��d�|tGRn���t=��)4f�S]o�QAI^i��/���ý��{$HhjF�'��p��쮬��s��+#�I�d>�͏H�	\h�-^��u�o����0�����zvq���9-�ӥղ��8�u���>S����`������0m8�*�%�<�,y��hM���*_��"��
_�7�E]�/��v,+�=�t�\ e�vgsh����F�1�(T�(�����%�b��L	^sOO�����ʕ|om�0d����5�yD���v(���G�����c�=��7�"i��=���i�T�&��PйN��?Mz,2�D*��z\3�Z1��.
�.��U��RT��ߟ��ʒ{*~M�z��aN��9�XSx�.;�Dz��n�§O��)�%`�"@�:fY��Db��S'ŷBž0O���4����W���P���|�ZŠa������^�I@~)u���͋��Z�� �Q�8�#J�ڌUV��I!�M�Z�_�*��h���M���3@05Ӄ�몯By4r���$_`*�̜��8�]�?��OO��|/��!b�cX�T�}��#��N�ds4�������.���d*K���Ǵ�Q$.|���*9�}\��?YfK�gY�H�JI%�]��t<��A�$�b/GZ�ҏP�Q���0�ZfN�2�z�E�I�	���ݫO�Nk�����$�� Q��(K��8�~��B�lA���U@�ăgw����ۮWE�6d��az��۠~� h���Putu�a���>k��Z]��eB�,��~�3������處�P���[*�OV"�w��%Λ0�I`���I���d�(AE�G����[ ԛ�co�U�~�#�r���{��f.{���_xM�WT�r>�)8I:�E0(^�[۸�ii�J���:��T#�
b�SUk�������%�Yq�G���x?���r��L�ӊ��WG��z3��&�Qژ��@I�J6�����Km��	�tb��h����+QC ���������&���
�,�E�-�e�V!b���#q���	�G�Q)�(��3rL������zJ���ߌ<	� ��ωSq���u��IF�԰�4E��E�j(J鉂^�%�I��vO�t*��W�,��A��T+�Н��T���ߡ��8ѓ���1�7C&��R��-V}��؇�sC��tW�b���iL���S�d�;�$%k��y.���VD_���@�P�x"���0�T$o}^�^ X�~M�Ӱ�/��*&�7�=ҽ�(���B��	�!;�o��Vg����s���y�i1Y9�fѰG��W����z��X^v�e%�"n��v-�c��	�\h�"���+v@�m�?�$F����UL^~�,��#YN�FD�O&x���w�-��y3�cw�_
.Ϣrg�a{/������i��WW�`�o��7��Gs�3�1�vD��Lf<#�������6�[�rW0~I
��W�����>�nБ�%���b�X�5�e���:�P+�ldnO'o�x��ߩlC�2���8�;�k���.y�Hbq���Jz^��Z�6ʀ@)U_:�$��-W<`(89�&>����B@z�����fN��Ԕ��������u�"_�z��I�:g���ݝ5׵�Ёp�iϏ��Я8�r�������I�7a�)
%s�Κ��X��\��][~�� �G|VV����C=�K\b�M��Xo>�ܲ�"��