��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D����gP�������������44��Pg��w�k�n�L�t�=�ʠ̲J�=�	�$tG�讧��p,��sC��Xu�_ S�	��mZK�qnu�*u"ǋ<�L*�2S���!��i�އh���
������)�=k��l��hx��I��} ���l��CaoK^G����F�HE���}�-���8���C��)�6v��q+���BɃ״��0�Ўl���Ax�`93Di�j�]��0x��uHo8ȁ�h�+���]�,L��uS��|�>5��9�8>�U̒ �|�o=���{�
'�[	��ԄgI.��Rs���Z�GݲB�_/h�_g�ˢGmYAa/E���,Ӥ`�΁b�d�@��+
��kz<ˤ(�w����0C݊��L87�C��������z��H�w��ڻJ�:>A��>I�B	�KW�-H��
 �ѶJ��;�\�16Ji�,�z}�:d�9E��_����Z���o-�[Ɯ��F$v�KG�%Z�:�oA4w�)[����:��z�X�o=B�e|�_2��ͰUSo����I#ظu��#x	oC}�v�%����KBU�2 p3 e�+�0ʝ��l�;$랉�A��t�h�?\�<��d"]���xuB�@3�{��e40/���GC��������ھΛ�HWR4��M�q��q��x�Gf�5�AW@{�-��LX�d��փ��Z�$�|�t��u�z(t�]7C�ua�Q�t��>l̘�9qaD���5:Ee��LsQ�����yEE����r�~eh�9ʋ�s���s'��{I���� ��]���±+���D�x��!��΀�����J����'V؎��`�������1�jvV�V9 �����+v�9����ٟ�/����I3d�D@��YT�ӵ���W�mD�x�&?2���c^L����+�����iP�-6���\��Z�HP�@�4��\<�Qe�gCa,���c�����+��Aq���
�*�prf��Pn,Aۄ�d"�� ���W�˙2�
T���8�&�����Gvã��
�t����{hA:ŽU�����>��J�<��8d|������ʻu%R�b���4�w��1�3QF��|d-ך��P���C1_ �=����kkH��RYb߿�c�����="���'��qf����V��D� K�d��=0��+x�i;	;���/R�Q�b1�ţO�Q����'�#�k����xTex�>�Ҕ�qХ�*\��^,�W������f�06�J�9'F���#,��I����2����M���m�RH �>�y�d+�ϫ���lӕ8h��o�S���GD�� f�]����6�Q�F�Q;��q����q�$��9l5�������o�Y����� ��,WPgyc��K7�3j�ဗ�_w�sFY�-[y��{WQFw��?ڬ�\WK�����$T������v�),��n�����Mu�o ��N\�p�ظ�@`�;3��<���Qٹ�7܁��ǫj���pU������0�*�Rs�2���na؛�-1�����aY%�EY�PW�Ms�.��%��'�=���d�����Z�4���y��4�+�بڤ��@��W�������L`#�a�>n�-�qo�U��-�-�1�؋���l�"���|����*�8gLd��e���3��A���#���go���e\��=&��YH1�.aNl���@/��ID�����> �p���͝�K��,�U��U�sp��E9�õ0l�˂�D�Ak%�F"�I>G]4 ��Z��tf���ke+�S�.y����N�J�ڒ����*�SI"t�W�q�����*�~0�Q1P�(:Q�j�*��¹��\E��r�c=�Ԁ��<�����~"ө�.�_*at��N�6B�1f^�.+Htj}@u>C����ȠZ�K\/	��橻�cl�r39@�-\"Y���(����,06c��S�crK1ިmY �q�h=��rK�ʆ6����c�Z���"��vL�p��D����D/p�����i�$��ϡ��s�Ժ�&�ᅴ2�J��b$A��@�ٽ�m��m���v��%*��A��}�aB�ISP��<PCU�ܽ�?W�`q�'V���ǋm�E�����]��:C^��+��f�� Xt�fSH��?Eg�a�N|��4ׂ�J?�P�X�">�P��S��%?�٬z��>�������m܍�-����a�f%�+1P݅۱F�E�}����ǭ�'c��T1�(g��mx��Lʄ���8$�g��C�VA$��a��r&�*Z ��ٗ�����^6�����"c��p�������Rk=&1f_X<bpG�����5��E-��^-��Qsڇ��gVʌ�`9ǳ�gr�l3�'2K&�i,����VR	���f8G����<ВF�R�#3|@�=�z~�^Wj�{�qCV�����Kqkʦ��)m�ȭ�=�-��cla����C�'f�%���w{�hȧ^�&�bu�G�e�޲M]XϞT� <V6���/�7ZWXD�'��+v�&J��'�,�l��-��̵> =A��]�����<0cŔ����C���7�(���F�_�[)�9���@�V#�h���;��a&�9<���ԆJz��aC|:"��C���M�ب�R�7��?%����	����{��	�$�Z�;�L�@��/S0`h�x�{p�����sv��6i}�����1`����j�w�1@C�Ǿ6,ԩ[��јT�ĖqAj�	3\~ջ�9�uHL����$+��4Sn{5�[����bY3�����L��G���%�g�N7��e��֠�	�@��S�������r����[,VY�i�A���v��v���ԕC\�v%?�0���`�뚖��p�z��Ԝ�!�(���R�� w�&�?4)>FM�z��}�ͪZ��,>_�D�/ʪ�R���	g�Qg�Q�T;�ɝ�۰��R�`�'0��zSD��F�����b�RB �=�[V�X_ԗۖċ�r�|I-S$��-��Q*h�=���)5v��X�m�^��K�y�� s��r�N;Ku2��ɒ��=�IO���������2<��=�.�n/���?yZ�e�@������+��sL�,nG������*�W�ud�B�z��)�������mP~�� N�]t�f /*�+�%+�r�Q�`n��\��׭������`��3�Jݙ�և�Zv��ש<X�_�FR~7JO��̖�/�ap�}bZ\hz�a��?�m�37� $࣏"�>6.4@��䕻�)O\��A�>惞H*�G7?�`�|���v1�������n)��"�$8t42�P=@�x��oB��5�W3���ʁ�|�\�մ��:�]9�B �NV�+�^�A��<��%�`T�`$� D���v_{*?��u4S64���4��l�}�`F�gKG��ʍ��'3�ŁMO-��v�/t6C��4���!��Tm�	�r#��Z=.x=&+�MJ��Ν��a�W��fp����L���l��x<�@T�K�D1���t��^�Ԛj�"Cci@V,���g���'d(�$r���ӵw�[�]�Z���NS���ĝQr,`��+�9G�Őg�J�uz\%�D`!����6�wb�R�Vf]�z��;�=�u��|��(EA�	sT��hd�ND+IE��q�|��4s���9`<��Y7�S <py �[0��J��;�?��ɷdzI�$�.�m��o!G��cL[w�D�ԣKS]�/���U:�����?PUWO}j#i_nN�\�Wt��{v�4P]Gs�@��&eNꢠ�ē��C��T��@�)��Wꕈn�z��6L�̬'�lv�sm�y��Y��ɉ��ւR�^=��������ȟJ'O	��'��j��ן��;�oMy�-� �!����(H�辚�:�?���D:�� zec/���׀�vb���s���oB��ߚC��ż�{�Iob.���Get���.������T5og�.�X�i�(�����/ԇ�S�74ϡο�夙d�)����4��Z������I
�˱O�5��`հ��!�
֔2�"���;�E�:���-����� �)�Zw�<y,/�K�*Zz'���ѣ��X9��8��D{�� �\C�RO�8�`�����yl�`s/xd��[}�șwdd ���?�u0�=��,B����'�F�J�!wTqе��B��g[{�" J��Y*,[Ó9��ɯ{:KU }Ʊ;�@I�ՙ@$�3����)ֹB���ã���\%��Q��Y�dd_�֋a}"D�.;P��s���j�cVH�.8��}�ʹ|1��N���S�1w�oN�4n�Zd��^���������D_�	�����p�}�B�k#b�a�.��iF�bK�����1���[=QT�?*c�
��K���Z���TQ��G�>����P+>�,����2뚸�\��O�p�����\mѫAzO��Q֬�T��	�z�#�ハ(���s�����P���;>=�u<w�@ڇ����:8ۀ�hY��j�c�m�e'�R�/�����#�3���^��[�@(ǉ��7X��G�Ğ 0���9��ϋ*�+�X�Ű��* }��jU��$:L
�z����M��Y �HCi}���i}\˪׏�,*�P��$��0,s8�l����:�K����M��t�$zdӧT�?�bA��
�%u��U�ǳ/�#x��&������8��^YΥv+�E�Q��15�E$ț3��/��$�(��[7c�����~�RH��|��]�e�����8��Dv�ebݡ���3Y�ܴDfšN��]��3D��m��^���d�3�XjV����N���{��uGN�	b@��m9���l_��eyfͻ�r��Y��#�e�B<=�D���{ý@���9N`��q=�����H��щ�	�B�yi5j��t��E̴Х��/9��p�,+�}JKN�&[A&��4ޘt���Z��O�H�C��o-����^J�%�'�)@u�q�Z��ek�t7�=��\�xg�c��%�@�O�ݢV�>��cJq�o�3�Kc1����7�u�#�By��05|?7�ǘ=��n�1C�d���ko�$�cDy<��9T��oe�R��vԞo��@M���˔`�j�<�̅	�]��sk�Z"$8��&�;ׁ�l��.'���#�^������pT�	�a<B��/ъa�����	"8F;��	J��76��IHs�w�vt�׺2nU<�?r�6�b3���a�3S1
z)Q�.M��r���g���s}���H?�f�ɡ(����Q
�֡�R�-\-��u���H|��6�L�~����м�Mg@yVN8����ХE�xMz�[�}��7~j���$�[���M�N<���L);�S+r�"W.�R��3�Q~������5�'g��Y���k�ߕ�d��:s�+؎0*Ep7�Qܿ��Vͽ^8P�W�*fzU�B"�2�dI�j���?�Q�0�k:�����_WH�=�8�
���<���f��a����O�*oÃLQF7�tBSL�U��獌�#�TW��tѯ$��n��K��e�T,�5��Ҝ�DC�4S�([��E�Tss)Ш,��`;����*�v�.�i��P�Wf'�<����,Ъ9_�5E��p�X�n�#����FҖ�}-���! ��Y+������3*����I������J]����W�WB�7�[aw�^��>� W��+����C]���4aD`ճÞ�i�2��Y"8`�zP�v1��
�\{��F_Մ��=5m�}a��y���O�A70\� �S
c�X����l�8�`y�*a�!4Ċ�x牚.���Q����e��u�u��ס��{u���O���x(&0�w��| ��Կؐ���md�oU��ݪ��D��m���o�����$8#N]����V���`w��\9sz�������TB.�>\6Xl� �sþe�4��9y�w���Ӵ�c�% ��)W�Øϴ�ʮ���i�P�"��i؛�CfW��?�fS�C�rO�>����oUr9;}Ԩ��3���{J���`@��?XǓ,�$���u�c#�6��4s�p���M��VrZ�������~8 <��7ȼ��[��+��䂏V�G�h7R��N�>X ��J��Xl�Б*-J��`~N�Jh;���x����I�PX���y3�'bΜ�WN�ׁ�I�V5�+z?=&�?D{q����{�]���N�f���[}XҪ=@� �|v7�1I5[*E ?������4`�������q��T��>y�Y��]�8� ��<�x�EX��B�n��J�P�:��Ͼ<��$���<6���u�1R�ȼ|�����rr\`��1��ӽ���}��s�c���Q�쓔;;����\a{J�
�<��P��B�JD���7R�$<�D��6���g������1�dBs���q�M2�t��?W������u^	Ij��U��%�\�;c�Iw�>������qJ��y��XMMp,7E�����(��-g�l(�Ɣs�4M}od�Wf�X���<\�/g�W�YG��/���0r�2��������1��Fb����<��\Wc���E~*ECb����X�J>��]t9�l�EYk���Nm!���7Xr�u�:չTU��ۈ�p�6I\fG�=����7��Ư��1"�Ӕ������ M�	�<�iC��yL�t��(�kat�ZR1�͛�_���w�������w�ҍ|����-q��X�{R%g��z����$��%^J�����-�� ��o�͟�ҝ8̌���W�3�$Iэe0��2�9�r9%��E�Z���!�
��}�󱩅�d߉��h��DB��m[/*��1�:m�t�!��pWZLB
�"#}pkl�?�_�Q���6�Ա`;x@��-�9�y$h3�EU@b���u��U�� �*��5�Rz"��Ӎ7����s ����
�%�8Mml�;�n�������x� W�=[/�9*��n��y�n8ےwI�gF���	a�ug�.S�&Z�/��Ň/&���D��r�w�w-����ã�-�gq{44\���/���C�s++��s���� �����U�K��\&5�B�A aDҺcx1���@���Y{��hV)+�-p�d��ґ��l�?�=���-���r� g5a�k _h�M��)N�y��y���!�r���!a��#��_�m ��3��n�?��p��-�n�O��[���C�����i�R�M�춞�}i$���7���] �*p�b+[��%�R���˗?��o*� @74�AE,�zL��Y��ڌ閃/��%>�OCúJ[�R�M�\�F^���NE������1�R[Z���*^yg+)\#��E,w��U��$����e#��6��)-z��R��vf�!���f����
ʤK� �w%� �{��3����dɣ�0rkT�9���	2a�h�e�
3�h���ە�/�-�� ��S:n|-D�6�Q�8R�bk�F�+�	���?\旳��H�����ۈ]*���4���z)�x񰠊��a0��Q�W5S<)�,�6F#eT��P;�=�6�g���UɴZ�.��tw��2�Y	q$]vnV�	� �l���@�:x��UJ�?���-�>Q�l�	\�掜w0(/L�2���F� E2S幀u_!C'J.�9^B�D�av�h{��(m$&�^T���:�UA	!����H��jX���3�Q�l�NW2�6a��J�� ��G�chG]�]�� T)���%���Z�d���9"��	!�9�C�]�5������YT��24���<��.3�D�:%̄+�՞`r�^'.p��I��S0��KbF,��b��볞�T�����Ɯ9(#[lQr򋸢Y#�1al�i���h�uw��Wsk3M�s�_�o�����v^��kUz�7FUXNu���� ����m���:�jQ����h]�K3���片P���跆sSoTB�N��c��(܋��igs�~q�r%���߰*��9:�`l��{��4"A_ERh|�b��]*�z�c�U��ӓr�U9}h���$�J59��7u#�'4�M���! ��0��L��)���Nhg���!�þ��>�n��Ga�N +���k�ᓡ��|���g���{����t�r��	$x�����hf!��k��%�<�L"��g�<)�ڹ�@�/.���F�x���7����5#�Y_�ه�����{�ʐ&9z�MxV�9]�xN#������G"�V�[)����K�,��U�Ⱦ"[
��`�0N�Elh��Y�%S�����}'j�0E�E�'7t8ϥ�US�3 U2�M.'ᒙ�
��-�����f��� О���h[z}
_~oTΙ�`���1^���r��z�gPƪ��P�����b.����12�v����DS��,��㘓V|�>���&pҲbt{�>�x���궨��Q�2Sdd�h`����ڂ]��	�^�S��B�:Oa�j��Ҳ?>?ޯ������a�M�ı�������,9�=(�EIW���91v�Hu+Uf[B0�|PQb�Y�K����.�����T^�����:��0����!Ų����A@9bh�	���Fõl �m1Q�tTR{�pz�����>���^�Ty� �l�.���`��[H[Y�EJ��1�V��3[��k����P0r�]�����������jbeX��.<���͞�M�:K��Ǐ�<���ܐhC���3��"��C�͔$����*Ԫ^��o�ptgx�.�j�#���̦��!"�e�Cqp�BM2����ԝ��_�{(��U^�$�3̩ T<
�����-��ǵ��Y!%�F����1��m�w��]��S݇��K;�,	�ƀ°��/���ZL-���]Ҏ � PBO& ��"�@4�-SB?7��Ғ�F����N�'����!���@�E�dr��QRH(G�|�xwmB� I[ԏU5�/�5m�]�g��^��g�@V-� y��	�Z����aO #�8���qP�<�O��$��}ߐT��z��C�D�t-ׂ�l&���W�I��Tk� �i8 ��K��>����|Uh� ul��CSp���r��/H̚��� �Y�k?,�Ҍ�s^��N�n���u��H|#���%l{�j��K��N�重`���wÆ�=��	iL��9_N_�JYk%E�5v̕V�����jeaf�0g�� �j�9�B���4��D�~�T���p*�j��"N���D���âH�U��j�a)�Iqo�t��8hJ=�h|��v��V��gU3�_�^ ���,�r]�eehz�s�W��OO ���Ϸ���g/ϧ���$��96��*i0O�0��PE�����H���tLT�	��I��[�n[�|�'��6rW
wkJ[��b����H���ᐢTܦ��t{uQ%�k�(X*g��3|�#&�_��(�ό���Հ8;��"IvP�A^��<#	�{>P!�����������>��ٖ�k��]�L�e^�Yv�|��?�@Еp�F�E�hcS���m�f��M����x9d}�fv0��aZ���)�Be�:��?��'r�{�E�j����zK��
�U�|-�='=Z��*2u��tE�߭��ɸW��{�Ѭe��R��!�6T�o҉N�h}�Vi'��S�z�'��O�/���� ��Zxlg#(.�d��b��f���B�_��W��9���m��� �G��n@DP`�A�U�l�	W|�)�t��)��1+�՘N�Ǚ{O���،e@�]Izv���6��9'����"�Nh��!-��n"�=2��n.�f)�� vHb=��1��gjbEP��;ٚ�I��R�q\��|��{�k�ϰ%2���u�M	lrU~·Z�K�v����ݶ~�3y�1��i��4V�V����b�l����h�Mq�� xi>P&�2�J��o2�����@aђk��e�؈��h�!~]�s���ݚ=O���{D1����6��H�m�Vm[A@y0h�x��=���}J��Q0��f�=S���_��}-Q1\����b���;rt�*�U��������N��=!�����̈́R�;��T`���FR��� ��N���J��Nx�D�G�,a\���F��j�6����X��\Z����}��U�e��)T�GB/�;͝Bp��wS9�_��t������jF97kW
8��f%�/3�w�U��z���Kξ�Ԓ��#����;�����Wb1ht1�g��q:��z�Z�5QDF��8oj�x���Y����t�س�׽�@�)o�^(�Z�`���k���? �k�u��nc��$�,B&�J��/;yR�ű���2��8ϟ�M�M�\�����JB�K:1N�y6Nv�������d�v��lq�vD`Ɛ0��U>���N��D鉽��]2�n"���5J+y_ޑ
����J����u�0���I��`Լ���e��XЌe:���Eeƹ:m�ԅ�sdS�&�|2����[b�X���XF�L��-���A�mh_���l1��,�����^:AOh��;��Ť���3�%W�������H�,L~�HӤ���RYL�v�M�WXo��;0�m+h�*1"��NM�;���eg{��s������[E-��1˃P�Zf)��v���Üd[��ܯ���R�ԚF�����T�]��1�6X�	q�� ���tL���/���g����ʖ@-B~�Bfſ�5�V9�[ ��Za�-�Uq� t4����R{|f�.2q硅�˳�D?�?�Γ%����/���/�@ k�I����a�u�e��ڹ�ݰ�#󮿙��~� w�<(���7��r�)1l[s�Ф}*��"<��T�J�; �!�5����D<j<kX�����N��T�G�jK{<�����>yA4�C-�	m��%��i�A�1�~��3��>s�B���T+|��^{�^�p1�m�bdֱ���0�%�����)�A	��:/R�:��E.H���?�$m��?;K�'>RN9$���W��p���l��(�:[���,���K�7�W�>~�?�ͭOܕ�E�hJG�&�7�r�����7��u0���m�ˤ0�����-Gׂ!��V`���^��M�E�-f������s	'�m'W�3A�!�� 3m�
��a��r�j��������
�W�E'yW̓ea,��󦃮���4�;PN�:vR��>Sh�c����C����3ݠ�K���@��Xz4`��r\s�et�'Q��b="!��+����>��O��/(�Pn�i��[lj2f�Ϳ��'�����(�S=����&��#��0V`Q�Z�����fF�y�^:��M�� bk���X��򂅅*��E�3�Q4��� n��lf�(K�?2�hr�� 	[����1L��!�K�Kky�i�uи��`}�,��\7p �X��3c��G�Ko6��ȸ��s��
]�`��͠O�9QJ_o��F��{v�SOB,�+G����L�Cx*T`��onW��2��x݉��`r��>4E�}��T�ZR�g�3�;^��NpZ�3�>d�f4�:�\���fnY�[��ș��gm��?��~�,Te����F�v���h��d
W��,Q[@?�?�]w���eʵ�=�p�8cU�쉸�I2��a��ڶB�@�5�.ǯy��r&�c:�О��Ԡ���"�[�Djs�6 �����:�N��v�^O9YKpBd��"��j_�Bن�z̼�P�M��BYJ��� ��]��cn�:����N�����x�wHV����_��hd2|��q)�=�$��$�\v)8A��$�I�S����^Ws�T�'����8Y�Ya�r��v�@_�4B4S�����ٮNE��i���V)�d(�v+>vM��7����|�N�N,��S��4T&X�d��$�A*����7�f�����5fHs�@/��Gw�D�y�껑�����]�^j�c��� U�-{L�h���uT�(`O��ز}U1�����2�*�v���/��,�d�Y�)�8<5i�"�H�ͭ����jxt~*^���n�O[��1�Q}[���cZ�P��hmz�IF�6��Kg�x|���Z@p�y��J�31�~]�Ϋ����r��4r�t�=��಩Җ3��MU_+��S{���m���� �������Θ<W�:g� ��L��rj)��G5m�}�O<�%;[�l��ڬ��
lf�"��d�`��Z���eț�ha�U��N"�Z�z��*ړ[�Ƞ
�D�t����\=Fv2������Hm�����b��Z5�B��¼��G����XJ����-��	s�u���a`���F�Vk��#�WT�����﹌O�y���Kח�ҍh�݀�5ƪa��M� WRh�
�_��� Ds
E�r`�L?��Jc��ӽ�$?I�+^��I%�e$�։��b4̫��)"�(��6��}��dZ(����"̀,�)vl���z��٭: ��ՊoW��0B�J5����@X(đr2CbENY�$Gy�b���j\�����%�V��2&'���p�{mP1���q��)��3��IA\���\u���W����.���z�dB����me�S*,�K4(�d�Y�W�ʥ���i2�+�C��/傰}6�=f��/����p��:\MȎ�Z
3#H�U��@W���,��ܺ�EƹJ�������1#�^�oO6wM�Ǭ���B�gh���!�>�7��Ľ��c��
ON���uRQ�d2����#"�;�f�ސ����#�t�ag�����$�	`�����/	L�����W�h��99��� ��Ь�-z��Q�7 �;F�`?K�yA��X�����u_�����{���#��������6֌�K�2��c����*ك�@�Դi�A�f�W����go���xQ�RQ�ʲ]jV�zZ���!��z�H|�SF�,����Q��Jx��,ҵW�/�(!tDt`O��R#G��ϲ�!7c2x�!k,b_�BTq����K`�Q5�d1�8�beGĬ SR��ɺHe�D�$<a���0����v��<��<֡G�َ�^�6!fd��� V�D���-%2�����s&�p8��%��J1�M�p���Z�}S�aK��2X��-��',/�,N�����~+G����ո���''}����%[%"J�Ф�yv�]�#Z��N]0w��q�9�%� P/ �ǭ�ynpJ�r����Ђ�����V�8>�D7S�����y.�<Am���>�O��Yұ�gkaa��.67���t��D�ϗ����s6���51���sG1=�M����-���0AF9�5�.o�T�}~�'���/�c��	p���{��f�`'��
ڈ��S���Z�0fZ�,'�࢓Zz�?$e Ä46�j(;5�ߴ0��6�(ϰ��"�0S�*q�I���������f��F't����j��߫�����6�x�����(�\0p�}��I��Fۿ �ݽ�ga����ǦƮ��<�x�	�qcSnwВ#g/��i,��,�M�~��>'S
�=�ǩ��p�O��b �w�~e��C�ցŇNWA6t�]��+\9���x�(U��D2�=�raX��,^,v��a�ϵ�+��C��z|�F�nvM65����V @�~��w��ӱ�q2}�Y�0Bʘ�*2+�ٹ�,Q,Η�,WHn#Z�Z�� ��lǕ�(��7��<$P�m1`^}�Ռ�,�h4�PL�z։�*Č���hi�>%i��8�J�N�!���Wa�\m�Q>��z��E���o�5$��|���!-"^���X�P�-(̗áUu�Z���ґQ{�c~~J ���BZ��&F���B�-Μʒ͒j��:�R�l��M=��k!>[M�JL�mZZc�EFc#��g�,3=�hx��Z
H���7���x`�w������m�I�o�*\3C���0=0��,��pۏבb��zĔ0k��욭��[���TY�:��~@�!D�A�����%(�K�����U]��C(����{�tZh��2�ۗ��}�.쳘�1�H�s�{��6:U��]�2�A�95��m[����0�S���S�4�� �@��5ʀ	9�6� �1<w_iC2b��~�Y��kJ�=k��������_��qZ@�ќ?���xǿ�0�3��hq��L�����5����s*!�h��[7�N5��V��۱�+��Oض�'�:���T�d�KT7������y��b@I6������g�-p3� �/~��l��{0�S��������*o3_u[J��Q��y����=��ʱ��TG���T����l���'�0��)>�ꄸ�5�����%�&��w�b
��C_��
<��GN�j���ͦv��R�3`I��ޕ�%�-�V���p6�� �1��i=��k+G>Lx�X܎�����0*����.`uD����>��<�ٍu�7�{�4�-E�So�����'�����ie@�ڹ�ݲ#����e7E�9j�s=K��+�bL���ǟ3f'e�<^�RY
�y�?����1�/y�c�@A.��S�#T�u�¡/n�?��v�sS�#g$'�1o)4^%�} ��5�f��矧���<�Z.k����3q����=����}9J�u��,��34�]xl����rQx��<��7��f��?{��T?�t�Sز�-�`�s{�ո¦��ʨ+k1ԗ�]�T"?�ߩtG;�8ݗ� \��}�����d����m�����<ˠ(R��1�''?b��I�~<x��6���.Qce �in���Wf?�>9ɵ�p�\�ә��W�f�}h�9�3����֬HY
QX%K	���
e[�t��_�Wy�����@5 �=dl\�M��_��D��1M��n����GS*��#Y����p��@���{Qw�;���F�<��wˢ�Jc�1���M�l�gZMzd�ve
B_ҖH��� PK��Z�48����݇o�#c��@��ʶ��/�LD*���ky9�N�S��������t�+RRT��Aʝzχ� f�S�m����	�-TT�,�?T@z������AH�EI����,2����3} ��T+F'&��P�w��A76��ϗLg��~@�g)۫8S�x��A���}$�p�К���Cf�śb7�����Ą|�lm�����Kv>�K�\����z:�������x"�+��@$"+�|n�RSu-Q��_7�}�H�{����;�< d߆�<s}>���ԼS��Q�3}FD�r9�c�/��z��!�=�5,�:��kjF'��K�<�=�(5� ��	�s��2+����~hf�<�j�����8��aA��q$��D�Ov��]�Ć&�.KcM��K�ݢ���S��{9�s������(v�$x�cO�;��2+0���X�B֪�_$�HD�7L��[=5��\�
{�k�6�y�r*�2K�V�2j=�3�	�j�.c�w�Zqk�W'X�k�a����s>e �b��l��?cJ��0�`� 0+G��(a��&�Īc�AG=��Կx(V���7(�&s�Vt�٤�/�3r�i��*Oa��%�#�<�Q�`��/F�Pߢ) u֞3�2��0Io1�>�I�0u�9��!|��<�Ɍs�v�o<X��W��ѐ��*�95��>@����}��� �9�.��Uv��G��B4�:��M�`������h���B�pɰx2\����P]����ڗ��IaM��(tBj锥����P!D6\n���G}��h]b�L�ǆ�`*$��z;�����g��D���:v=6/:\v&M�"���U[�_UPE5�N�tU[v��Ǜ$_f���ߊv�R1� AjX:ڔ�d����~��Y�y�#�3z Y�s����$�����o�r��zY��,� �k����p}�r`�)!pc>�'�c�U�;hJ	�k�y,��H2������-֤SZ���]�6}��@�iKp�\����ԶY��(�g8�lk�Fu`�]dʟ���ds�����슳��%/J�vU�q�R׺�a+yr����-��.����W'����L~��뮏��ٗ
������H�ԸTK�J�s�J��������ؙk�3�{�(n�L��[]@:��:�R}����~\�'}��il�r�y/�F�o��S�E�]�"�M;W��}�4H0�9����>�6;t�9�� ({��/uF�a�'�n����v@��D��A|�S��C�8<���R��ә��5,�J�l�^w�̓Z� �ܠO���n�X	��Fu駿�rS����⿕>[��"͜�QT]m7�ļ��d�`-�W�:N�ԣ��_�4��1#W��NY�U��X2�� F�R���S��i��ޒP2���'��Ib�$@���9���Q���/#?���-Gֻ˾�����(�U��)�|;�\�����̺�,�E-�������O��7/�wSp�f���w�m�=E���6P2�HO�����f���}�n�C���F�^���Ra���J�j�o���e�W�d�4�9'�/��`?g��[[�LxX���uݤ��fO�j�㾷\�Գ��������B��_��#i��]#��/|�ր�3\զp�j������,��*�%�;w�fM+����%n��<?��Є�zR�b�2
�+�~�!����D��縨��sB������躁3%���4��
C&'[C���!2I�<	���0]q�Z��O�Ng\@���4�o�N��گ[�a�@bkS�N�`	��<��)�ip�tn܎���(��z��%����4��w��x"u����T@���%7ZY�Ԥ���;r̺�f�1p\��_���>4�$'x D2!���;\�`KG�b��qf9�ߣbv�
S�B��@	=0�*�����p~@�ۊ��	u�~�����}Tټ;�X�
>�o�r!4������̽��,F5��R6�� p��4*��X�t��G���J�e@��@�۬%F�ZpaC�P01��K�
�H`�A�|�a���'�����q,8��RnՅݍwwD| �oXe�ƞp��6�X �0��������M&�8 %8��95 r󪽶���}�x�2���g���XWd�c$��q���ԫt�­���S}�ѥ��
�|�YE$�Ď��0p`B5�G�M��#���3/��)!b
,�޽�;�Ή�X�e�'�{RΦ���}��O�9S��ņ*���f�L��Rh���J���H�tAd���r)�%�d@L#2�$�9Pf�1�:�w�A�	�	��c١��Ʃeh�U�>�Wr<�:hu"Ӯ�+`���։�F�x�ua�z	�tB/ӭ�
�y�1譸��b���S�~���V�H�O���r��$ �(�	i�+�,�R.Ր�_<Ԭ�W��N�ìܳ9Ƒr=����62��N8ڿ7� %����n|�jh�36��zJE��P�塪}L��ڵŲz6�~����{��f#�R�$�G�$�d�P�b�%��IL�Zw�c��b�9�<�2^m�i:��hԆw&���]���6j3��X�+�Q|v=6a��ň���/���`و����qs{����>���PΫ��b;�
�fT�V����"F���n�GR.�Li�"j'��w�p��?����G�Y-�WS�2�'?�96N��fP@��W��)>�G�vK4=Q�0�*��Z��/vW�%��I�����V��2�%>�Q���ݿ�Ӡ;��PܿIY�uSO�t�Hƻ�	����2�����(�Z&�%m�6�M϶�h"ಂI	�����=t�7���)�J!$]<���{���T�X���kl��NM�Zk��<�.���ł���}�@�{m�%]x�ۅ���s{���Hʍh��{]�Fa����1h
�L5N����{��JK�#e �qV#㜆��*�zSa, �"DݔO�Cv�^JR"3U��I~Ω�ą��b��z��jq�u�lV �Nk*��?8N��������'р����t��
���X��y�����t��w�+*SQ�+6A��Z1�T�a�Fw��:A4��N�v� �'��T/@Y��e�D���������$۔TBN�� fq��ռ2�D2*&^3��J���Y�p�z)��Z��(�;U���x�&�ȟLܓ�U�}_!�;�DZb���vk����:OX��]O~�����\���5l];׍�	Q5������K!"��tZr�L���4���A�b�����z����FO� ��H-�� �xqs|*�*!�2��]U��R�	�K�Ue{�����Bv�@��qcg��_P�[��n�x��-sJ�o{�����ġ��zy(8��T� `F�w��Y���/��R3��<|c��L�ʹ��bը2��V��1*���J|Y�����#�h߅��`�o�,�Po��� ��ێ��@`�H.���E��Y�� ��	��*?��t��r�&�u&P*Y(�b`Gk{V%�c�Z��&�;���LTVL��aJGiWM���� �S/J��,�Y�(+�l .lG�,�2
����Z�CYr6�]&.�>7(Q(7�MR�H��3�f u���:qj��aۍ׈��n\�����2��:���-��D�>�>ג �탒A��)��	�׻�r6�F���n�d�Cm\��V{��:�8G�o̊��\�q²`�Eq��iҁx�����2�?�w�(��k`Z�~}iW'5��L���~rs��7(�\��o�̫���������56���U�x|Zl��"+o��Qk�}ܦcc�Ђ��㞡B�_�xW7>����N���n�/�=���s��=���Pd�ZzF�T�뮹.�C�[]05p���+�Yf�mvIV���!v[�wrM��({���p�d�lc��X�4�b��ή:�B����@��f�7l�� ������TTO|K��Zy�� PYwLn�p�'���E�Z��gǺ-�-@�t�P"{[���̞�}��_�rd8���V�G�@IQ� #�rcm*e���� to?�|ƈ�\��TJ�9^�0��q���Ň��� �â+����I���{��Ɣ�;���y-hv�t���cE����|���,B8������fY#�B��� �C��<U ��Z�eZQmUD0���Z�\�k�-�K�k�����ܧ�~rN�9��҂9$��S��Aʈ�߷�ί c�w�����L�HO���Ρ�����>���?aD�����Z`W�e_K�GQ�B��z�6� :P/����q��g0�%7ߪ F���+\���i4D�(��dN�	��3R��h˷t��mIg��?���t�=N�ٿ�묞���PC�@���p]AX�H�a"���!ѹ6\�G�cY�#�C�D��U��G�pF�n�
X;�����m6���0*����|l����Pb�>�7O�Pu�0�S_�oT�cLu��{Ŧ�M@�HPҩ���d���?��d�)����<���{���e��sP@��B�{���!+��|2 _P/m�����Β��C�?��Sb�V���	���\�!t�n�o྿Z�#I9%ll)=�[ۖI�k�FdN`)*�Tf�O�})x�(Pp9� ˶g��i`2�C�� �=r�˞�O9�3B+!�3��9�.'�C+ �Ӝ6��k0N�w{�� m8pwNzK�` Q�)�b���=$�]݅ƨA�E=�ko�Ņg&�w�5�,� ��y5Ac\��mg�"�_�6Q����[-�i�#o9d�l�G�]�qT5�	���#A<nk�I���8[ �LS�z{�����r��y�P�����.b����_��w_pt2n�s�@ΩB�T)�rgF�A�- H�����i�Q�*�Uz���Z�0RY�ɐQNx}K�x\ж=g�[� #2�KMo�Vs��U����f���+f�*d��3�Z���*��B)���w���6ƻLg�q?� ia�մ9�Ɩ"���N�DokH�{+�in�D}!�۞߹	����nZ�Q�D<��.�CI��s�K��� �|���y��D�#w���[T�	Ez@�Yc�	X3l��G�!�l|�q�+�v�����k��?6U0�����H��������\��F���5t�0w/�D@�95���Z�if���:O2\D���L�`�f�&`A����<�a��}��QH=��a5/��;f��I4O�0\QJ��1t����N�zD��X�����ˎ��ŕ��-zE*���������ۼ��y����ڶ�p��4�g�Q�4�:��6�E�F�Ӆ�po�N��m�L(Ӭ�*���Yx���#7�Z�ҫ�7&R�?��O��^�
J?;5`C���Ù�q$j^��j�O�Q %�;�q�gD�E�w6��^g�(`�h]��)%/����q\����S���Z����c�2)����3:���W�d�F�+t��޵�$�;'Y��7"A)�-ݗ��X&�L��C�}T��A��$��,�e�3[�3�ַ�k�_�����_`aH��{�_Ն�;O��J��e�C@j�䆋x����Оg��8WRzi6��g�7"�j�Dx�]>�0�*��-��4?X@��{��泡,ō�{�Ο�1��t���X��$o��ͩՖ�_��ҮR]�t^^�Q�J,�����T���:���(=�&e��f�v�ɮ�\DxG~#��`��`�S- �zZf��ֿz���f��-gSR��y�>S�2EC��^�� ���(�B,�Z���9eiښ��Bu�s����nۏ���M�Jn;�a>�ݖ����ȃ0p�`�eD�xR�:J����aH�h�i�M��Z��۷ؚ�����QF���'�y<@P5�ѿ#b__��bp�h�x��/y	_p���p�l����Q������|�ԟW�w7~���m��֘�� L��dkST�������� 6�ЀmQG��`%�<!Kp]�t�:m�IZSV�\���J��"z~5{Ķ�-�b��s��E��V������œ�~�b;�RH��?��\@^1j�`C�|��E���� �]�C�K��F�B�ŗ��0��z��-�涁�<��S}��tX��1�q�|�
S���a{��M�"-g"ωPi��8����,F#(f��tf�_��a���u�)�F49�U��7u�
�FI;��	I,�������.ԕ!� ���(C��Z,�(��&.D*�q�ب�����gz�kx}]nk�o�(��e� �E�oeYjW9�%��eβ�¦w���2�Z� ���`�8�wB��
�J�$G\8�=oB��^ ��0�� 'N�����`4.l��?�:�H4��F>�a;XZ{�Ɋ`oGU�/����!g[�3��2��qw�9��3)qif�*�Ǌ ��p@�o5���P՟S�;~H�0����<���O�l��h����RN!^�ݽ�v���3��Lv�=��������E�Ě���F.��
�^|����$OyFK���d�sN���R�]�/"�����r4"�7����?�e� ���=�[����V��fpR0Gyi&4��,^wۺ*pL�