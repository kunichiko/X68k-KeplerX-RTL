��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#x��,��bZX�y�l�ob�ǡw&��2���<��n��\#�i+ ��ޯ0�F�VUW�J�'�v~��7� P~Cl/�MXP��>�g�!�iG1q��� �j9�����/�<�9ь��t7)�<�lvg�fg���w@��>>\y�͐�e�3��������t�7+�ࣵw�����	|C{�"r�U�(�tj!����a1Cϩ���J�s& ��@p
��Ѱ��@�2��d���{3nC�H�2��7~��wj<�v(��r£���
R}�����V��yTASt׷��l	�E��a/���/)�g tV�"��S����Ҍ�z�*z���Th�	Ʃ>K_�ϧT���'%IY����ܢ7�p@�u�I��V��D1�KZ�'��h�\6?��AH�Nr�P_T���Y�Qd�tM�\-j�"0e�Y��V�Rr�=���Q�l@��t�}��GZu�oŃ���ך�j�&"��r5K:=��S�\���P%���>[�5��"?�.x6Z�`�q~�9�l�zŎ�I���>�L�&��˷�g.��ht�#}d� ���&[��q�93$q�>-U�����q�q���M5u2�^�1v=8+d�k��;!v�x!�Y��lx����N�徂��Z��r`�/�-���;�����DO�w���עV3����+�Ly娂��D}�:i˝2��Ӓ�!�I��՛l!z�~�u���P�3%�V���a^�ۋZ3[g��\�����lK-�H���[��w��D����z>H�%��^E�Ca=-�r$mȒ�������0���4�O�na�B�81*�ϣ��k�ɔ3��z_o P���L�:�MF��ݦ�_cK�H��8Ȝ�{��T|c3��E�k��_��]����|)r�l�H,�&_�O��-n6���&��D]��G.�0!�;>�f.�"k���۰�Et�p�Gi�5ITiY��sP`�_�c��<I�P�Y���]@P�Xȗ!8Kkͧ��H@"C����w�����j�HZH�Ժ��ɘf3��|��t�ի;�W)Q�T*Փ��J�w��5,��A��,�F����	����"��SjS��0�As�Q^;� �+�q�o��{�a�gڦ�̯_\��7���se�=�.ĉ�V����2}�h1F��eiܣ�)F[=�r�;NQH d�T )�Jo�md
���h:���}��B	z�Xhd"�z������-Ҩ�9Ebqf<���67<���7&�;�(-��h���#ׯ�Sľ%�r��B�&���(��:5�u�v����O�7�@3g���<Y�ts�s����v`�g���<��3�2�D�<@5�-������#%��j=��9������Dj�J<:;��ȭq%��@������k-�,���[J��{�ٞ�ʩ��p.nhr���z	�1��S�ڍ��>�$�Y+�iA�$R�5�|q�q� Q*��?�i�CS��<�ȼ����ǲ�Aއ��u��,f.���Ѻl�P��\l���˂�T��� Nc�:��&B(b��>,M� &i�P����D'�|[	����Ui=�V�KW�E_y���t#��x!��A vZJ�?� �m��%US�,W�
�=�D���1 �3�#�����V5��>R�������8X�z��`��eT���c��mm+�E��	���s{Ei���+2ж�M.��v��q�u-ElY8�ܙ���S@��(�nՙ,IH�9I�ȴ�2��}8��ǰüv� ��g!�]I���~�k�>آS2�����n_	zd8�A[�mh�\/�"c���[,2�P��� ��/W�=G���%kZ�i)�'1�A+��ƃJ7��h��stn�I�c�+�P �2�N��sî���M�k	/SB����.���l�8�,�$4�\�rZ)�{�5wT�e���SZ��]7ھ)��R�j]|'�CI��:�5�C{�ɨ�8:�?�F�=��p$�����ULQ��T�攚�ME��H�a�W���f����>3�*Rnx�V��+�������N��%�B]�����a�1��ʪǲ�w�*�&w�y�d�c�	��(T9�x��6IJ�Ư���Р�ɩ�I�D+K$�oC�+��CEb��#z�.��u���U���E�B�cp�5����0a:B�n�4�d�A�2�I�%O(�CK�x�eҙ�%ՠ��e�K���iG��<��ҋ8�Lnޢ���Xsor�>�a�����ok�:�t{n�q<�<V'�JZd[ʫ:�w�Fq�;e�H�Ո���(����iy#Y�G��$������h��εVU�_����`<��=��ex�'BK}��g�B�D�ZdkP [x�H7���^<�*�[�=Lu����
����ry)���"oه�wSM#9Li�	�0]&��:z��i��� �qŘ���Gyj',��t~�%o��yd���$I�Ϟ2�)�xo:tl��))p��e�AU�P1��ܕQP�yD���LZ(j�Z}ͦ����0����V�}�^h�A��~�.����>��oeD������Y*iEf��1�̬,�徲�R[�Mz����Z��"�"�v��|m8:/�Uև���)ܦ@�®�(������^��+
�����V��儛��m!w�]E��25�%��e��t���x�P��g���A�����Gl��h%P�,��7�n�%��z3�Q�B�N���K�a���%A��3I����oԑ7M�=E�ƛz:�Azo�.��w'))�4p��0�E�p�"��u�>m#
�lE��r�o�m�P���H� 	A�~9���zV�,��M�d��6�GM��Kii�-'S���X`�00y���87{�ևb1�{��'����!��Ɂs�P�$>*�ݿ�{��l�-�F-e�7P��Nm�*��D�ì�O�Sc�x��U^pzϷ'�z�z���ݼ�>q���I�Y;�?�KX7�ʤ�d�IyR&9���|	����̜������R����KV	+��H��￾�A�#��l�ou��0�_�d�[�����"A~���
J!E�۽,q�l���>G{���%���3Ս�FY�p��)�v��qY��^G#�:�z��'ҞA����Ӓ@
�*�_���
�l#ԟ��}���^u l�r��m}U¡�T�Y�}3���!���&�)!����gۿ�M�z?�K�kB�n���fۗ��(��l6߲���(�6dm�ӊ(V̛.�k��\/6�!�ʸ��3y���"G�ͫ=x�_����\�߱4����6��/ 2߉�!r��,LӠ�y���6�ƅ�*
=<
����1��17|���/���H�@L���m�2TRR�����/��.2��&g�	V:)3���ص��:zI��2�׳���(���f���W����d��nKBMx��&&�Q�&� t�#7A��l�?L�E+�������C�=ܲ%�'� 6�hhe�n��Ԓ����
���h�xZ���<{faoB2�S_��$]
����Z8����L���2��h��������{�>x��* �O�s�?r�V<����
�;��e�P��<���J��6H��#{qB�a"/���O�gX=�y��o�=w��������
��r���XIhk{��Vda���d���@��O�$�Ԃ�O�T�ŏȟ����q�W��ȃ쐒�|M�����P���:�Ll��B�\'^ ��M�" �(;=ܘw�g0�1��#yt�?��9�Z|���|�̂�-�cDN�-ё�g���$r�!=:�� ���Ǫ�ؽZ�5s�B�~�jJ�>��6�a��%���I�=�1�����I�23|i!n\�b�#�
q�CR���{Y0�����~�	�]�<��7YIA@M��w�>����CRB����.��pC�y�Q�N�����	<!��xU�75�|2�z!��o߰.p>/=Lbzm��WZ#���s�yGcxF�,� Y�ܝ�u�	��c�*�2h�E�=��I&���5�b���ܳ�Q�pe�V:����@N��}���^]=��6`w����Τ�5�8p~�k��9�SJ��'�K_���xi�Q�F��W��I�!ʊr�m�Ki��b��bO^H��z�:�� gB�%B��0|�R���뫪ݟt��6ťIl�1~s�� (������.����2g}_���%GX��gV���ð��G