��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��5�������B���8���"���FE�Ҧ�@�Q\_������C]���5��1)2���� hڻu1ǯ�C�ƾ���kT��_W�p.=�@�0�l!�\�F��'����e�4�Cd�����Q����ǒܝv�D�w�l�!��V��<�1�U��Տ!E��!D�6�4O}=E�t�ՙY���#c��$TS��.�4`1f�ZG%�?4�x���<�!7��1��&��H,�Q~�&t
�d��M�p\�|=
F�oބ=� ����~Wx��5G5*ڥV�	����J������<�k�	�]q/�\U��;�h���y� ��`��1����ޒ��ſ�U����}���-V�-�̫��e!�r(���[�!5GM��A�ٯs%�Ӻ"�z:�r�2$�n���A�F���4ù���A��P�m�M�>C�F�����<A�>9"�jT�`�4pR�Wk$������,h}f
f�6��ﰔp^��?�|��QK5���+6� Dr������ޜ�h�_�V\ڊ��O;Z�>����B�dء���?�]�I?saZ��$���Gފ7<�{��Ø3eu(V����c]���O%L��kI\@<uj2����&W�2Or3j���^_����䧂+����/��? <�΄k�${*�����%�;��'AO��~vߐ}h5��)�M,�<�ܢ�un'�Fw���,���d���Ǐ���@���[͵cI���p�A#�������8�Uo���P�֯�Ri�N�JC�v��7�{弡�~�O��V��ۦ4�9����k-��b������Š�J�b�������6w�޷d�d����<^ ]_ƙ�	8s�Xc��e��>ێ�"W8*�L	�c3
�N����'�nK��EB�bl�)5v�Z( �i	�+;��>��x$P��)�=E���(�B�"b<�BqX��ʼ���ydA��}� �v����Ct=��Ad�:]|ϯO���Wwv�u�y���wpTOp5�4j���S�*�׶�C~�D����OZ�w8���ZP�ل��;���8�^����)d������ʿ�w��"P�J��tFC�$J��Xl��]]6��?5����?�ڎ���zO��aZ��?��С�²��X���G=�K�R��=�3��w��W9
��͛]J�h�G3�5����q��r��0T3����/�Wy�uD/y��A�:O��
?7zh�1��i'۴���R��v;';��6,l����.� ��*�(�^j����ں�ԩȦ�6���`:����. d�R�M�N���
hP�{VM���n@S��E#T�45B�[����a����lCݠז�A��	��F�q�E��)�n��
��D�r��/���ܫ��"���;�b��7b.���(N�b~�MU�������r�}�δ}]�n/�@k2X�.3:�"Tk��r2$M���� I��X�l�5��\��ݔ�]���Z��3c�@l�۸4�޷���H���h��`�@`W�V�gU�����nN�}�d�X��j��@��=,��Ml�f���	��&�Y�y�5(*�t�l��	[�G]y�e	�߷昘q��&��3��U	'���lJ郙����Ok��2�[�C"qhN�}k<��w�z�)"�Ϣe�d�ȧ���0��o)���)��ї�x�L���7�4�ϥ�#0�����	Δ���t{��(�I�148t��v���8�Tºj��Sx��I�_N4GU~���'!���,�O�5�p}~k�0��$N=ǲ��WG����חf�����A_�N��[?	Zh���	�����i�k/$K�H�$���Neg���x�4�6�8':�x����dQЮ\p����6�����Ґ�L�&_�:|�<:��9�ZX��)"��w���ق���]ybK��[Lm��.��}-�=b�|j��.{�̜������(Y���=<W5�	�C5Mu�S"��8�ˠ�����z�;n�+�r�0���W{�������\���Ҍ@���E��kJ���I���S�Q�k[���#^������Xp���'��X�ұ�TY%|ţ{�gG�}Mr�*
��)o�����4�dr�K���W-��EJ�]�}�\�a�O���O�y`�y#rB��H/G:���S9��*ͫ�c�6|�j|������aغ ���Izʬ�)_�����ot�8ﰵ��g����yut���^-%��R�{'��YH:eMQx d���F4����7��$�ƥb���ot��mEG�A�^�	��C��K	�c�=v��0	����� ���dK��IL�Q��lT,Y��~���6U� Ef�W���u�t���rA�܌���+I�d���`���H�Y0�|a�9�P$�?�� ���x���
��.t素=��Ҥ ���{���e�(�M��Y��;ΰ$�>��M���#M�S��F�={�����N�8a��¨����tY�j��$=� �������_ms��J��p���T�qoY�����n��G������^��@ݝ�tԽ�Fy��H1��$�v�KlA_zpT���#e.�qJ�=y�v?J.����z�#/aC�U�vq̴�ޛ..J;�bd�_�(@.����p����c/|�Cb9z��1kO�/������ӧ��"/�ĺb��ƗśvK�}��3��hT��¾��*�Ux^;���!"��o�!���>�씣�>S��ʉ�'�匝[Jߡ@WAn+$��� $����hy�RG�@:�!�J�~�ԃ�WoƔʌ��_��O֊�T�Ji�;G;%U򢷭T`��d�{q�X���ր�L��z��Zo�19��y34���P�I���Չ�f�D���?Z��C���6g��;�F"�ԹgN�G
Ӆ�����[Sۏm�|���e�<CA�ip\�� g���S��b%���-G�`�59��T������p~��%�bو����|�H�-�Mbjw?�����)	����곳���z$��`r�rW�aZh_�M�$����17	��[U�w;oW��5ɧ�����O%E�<۰�V�j�Lr��SK�w��b�2ab�-�	����U��:EvT� ��*����}�u\I�Ġr��
WM�+�Ga���ʝ{�-] �#a�P�8?	�z�#�̣�@Z�x�;&�#��t_�d��9�lB�¹t�[g3�y-��^��ضH�sL��}����D@s���n<1���+���r�)WVS
�X�W^�{��w;�f�/�z�̢3�����ĔX�C���h�G��E�zKjk|�bă�� � �
�� �vU���ɛ�ү�)_�?b�ͭz��Y۽����	p9T��Ú6�Rw�k����G%^18*ј�� �k\�&����{N��/������d�@��vɇ�Yڇ75��7 ����j|!ؚQ;�{ׄԳj�[��e�-ߍM���Y�6�_6����~e�߼sS��{p�`,!��w";�R>e���nb�>&��b�3������n�3�6���i�d�7�����VAk��GX۵>S� ��bk`�[���ݪ�k��*�����v�$�����D9pM��k��)�<��֝��������g0L'�	������TI':��
k������I�L�B����3�Ã�+eL�?s�M���Td��v���M�Ɠ!^�=R��&G\�I$Y�I1�ީ���Bb�=L���4#�������6�v����@��b'gT=cVs}�f>/�о� u �(P�QB3Q��9+h����%�����	u?z�`@O�AS
�*L��_��l[>���_��R\;w�C�N�$7�k���Y־D?pOH�N��D%
��W��r�	��6l�K�b����!�G���f���x��.��c��E�k�Q>Ņ�7�.Ȉ���h�Q)�!�[E�Q�G�4�5+M�*���:�^�ֲ���8��$�����3����e2���٣ ����H@;ꫢ̩�B�u��A&袻ҽЋ����C�Ox�Y��4m|�gRY]��F���7pzP�ʭ��=�^��'��{T�n�+��02����Xi`\5����ь2Մ�tj$�A˨���N6�f6�wփ x���B�|�L� �2���ɒS?u�E&%Kԙ+q����7��L��.��z��:�z/��-�[�b�j�=}��.N�Hj �mI�(�U�@�3���~x����V�C���`Y�*�J��X� ��v��K���"q�K>�����qA�)�I�[�tg�d�R��Ӗ�FL!�թ�`��+���cѠ�ae��C�K��}���L��L`#������$C,�G��6�S�շ�4�L�<�e[����O����������f��'?Ѡ��v@���\h8rJ}����� b�a����D7�#!���*��ZD�� �n��S����������!��U�^�N�4�)�6��]���V�����Q^w��<�v�ޑ�/f&�Wp~뗟�h҂��P���3{ǃ&$��8�G"'a����"�P�^56�	���B���ɴ��[Կ��kh�
K���A��:��~Sg��a.�s�!�`~��r~����4��ݷ���e�G��ؘ��%���7�P�#K�6�RGM�J�qi��[�K�Y���Uu���ϛ�h��S��Ĵ���4|�"��D��(����k���
���4�+�R?ym��D��Z��J,�JCO̜7|Pw���%�Pi�������-gC� φ�k�C��W��ҷ1�/���Q�q����êz�0`�5��{��,�vlj_�R8�O1Nw`��;��\#NK��-a�l����w�����8�Rg�M�O��S��A�\�XG�==z��Y��;jPi@��s'��1��-?�`���Q	����"͈��!�V!�?�h �}������J���!�H(@���gV�A*��,�妄���n����*��j���l��b?�§#��m3o5&���Qz���Q��J��99�]jkG}n�S>[4���YN��T�%�n������u�=Hs�iu��8�*��P$���A֛�)������g��u�� w����\$� `�F�a�ew}�_��u�y���@󈬋��wt�<���@e"`rb�*����KEx��tn����u-#vp�����n��-���Z�����wJ��Ry���ˮ�����_}A�1_��;����\�����4x(�]N��|���e��3(���zYK[�/�����b�^}A�?�~�9*��Ls-����t�����[�L�傚U}}(��닉�]y�9�\�!0�,�RVq�us��>�&Pڼ9�cz�B@�L3p[��2?UR9�D�I�0�Τ6DH���
c�(���A��Q�$7���j�(�fO"�������
��g�)��O�1 6mަ�,H�t|cl,3���(�+����.<�����r
�k��҉c�/1��N��|�f@�ɐ��K!��j05�Q��m��f�v���a6��Rg��"�!�� �Y����M�6Gۜ���>\1C�`łt#L��^��a����C�"�F�G�~�H ����i>�>���F�1�ţ�(C�B�/�=�'�S��C�P�%��u��Z1{!���:����aɿ��e�u��Z���ZrB6-� Л�o��J{�r{�	8��4R�[/�]	j��{^�n�H��k�NQP�+u�~
 ����a��%{mє<� �[d0����Q��W��_!����U֙�����Wh\���iZ�����~x)q���T[�IWH����}=�֯������$d��g�<���|^s�4�����F���B৾[z�
� l>2��	�.��IP��x�2H
Л �)�vq�0��
�U)�YkO���冏6w�,s�͔-�!~�EëM]��j̼" Ǌ��A��) �A����������`��э���{ !��Z�Co?��$�óS�4|j�ll}\�����E�U�q��N�p�g�{6���P3U�-�s��v��^LQ$�Z;���E��E�a{�CB-��|JEc( �����  @WN"���6�&^���P9?a��Z+O�,��UMRk'}Y	��	��츕\cJ��;��'H% �?�y��AdЎ�Z^��/���<�kpv�{չ��#����$2��'0A�V)(Q.��S<s�S�}�;�OBfws�;�F���A͈�
tw�q�57�H]4����������A���Ĩ�R<�z��bz�+��/�T��-��V}�c��j�|{�����>�	]�z"Ḣ�I���k|���5	G��ف\��Eˮ��A� .~��#!O�cCf��O�Dc��L���ᣠ�3s���f産T��Ú����X�9��W����oX}���x�PS�b��8��6�y+n|;"o?�����P�M>{j0�n��n�U7�	�����u44��g�w��O�gY��R��Gt��r����1:�N�2bE�\��P��H��*�g�ĥW���^��m�|YҭJ��J��ȿr1�@܉���r�����mV*ؿ����,��4�ayTJ�~̧u�ɤ�XG?���:��d_��J�W<	� ���|QK��_}��i>�0�����׏#����D
��672B�|k\�V����I��з��cU��?�Q\������M�GafF���hѣcz��k�SmC� ���j|4�K�[�d��Y��!G3ܒa��9�7���;T<{į�l�!� �!*�׌�������m}� �{Ƙ�t΍`Fʅn3Y�C+N��Ί�s�c>�2�40�e1�L���5F�$A��e��I���ۉmU��}����P5T����oH7�m��3@�J�z邗�/v��\���x����+3nVX��Z�b�l����2�)L�m2���`�x�ЛF�% �-_�(yw$a�{(q4L)�����w�E~�Jq��j_� R�DE�M�*.?/M���L5"p&�$)���b��3}�<�" �Z�ux���>m=bO.d�t�BB����0/���~�����(nA����Լ���u�y�X��g�%L���~؆v=�HG76ϪuWz�����Ĥ�0��4U���{���G�/��lQF`@��Uƣ���%5w\���53��0Zh~P���s���W��jt��A-�Ն�^�`$�-{�l�QZ�ekn��0��?G�}@$案��.���D�SpOJ'��}�׆m����W�?9		]�O��q�~˗x��#&���%����?��k���J�w1���pw6�rN����V���Yh����Jryb=L�A��#jw��=%�dK�q9(�<�'�wo�h����%\KT=e��-,5