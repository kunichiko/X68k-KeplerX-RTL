��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D����gP�������������44��Pg��w�k�n�L�t�=�ʠ̲J�=�	�$tG�讧��p,��sC��Xu�_ S�	��mZK�qnu�*u"ǋ<�L*�2S���!��i�އh���
������)�=k��l��hx��I��} ���l��CaoK^G����F�HE���}�-���8���C��)�6v��q+���BɃ״��0�Ўl���Ax�`93Di�j�]��0x��uHo8ȁ�h�+���]�,L��uS��|�>5��9�8>�U̒ �|�o=���{�
'�[	��ԄgI.��Rs���Z�GݲB�_/h�_g�ˢGmYAa/E���,Ӥ`�΁b�d�@��+
��kz<ˤ(�w����0C݊��L87�C��������z��H�w��ڻJ�:>A��>I�B	�KW�-H��
 �ѶJ��;�\�16Ji�,�z}�:d�9E��_����Z���o-�[Ɯ��F$v�KG�%Z�:�oA4w�)[����:��z�X�o=B�e|�_2��ͰUSo����I#ظu��#x	oC}�v�%����KBU�2 p3 e�+�0ʝ��l�;$랉�A��t�h�?\�<��d"]���xuB�@3�{��e40/���GC��������ھΛ�HWR4��M�q��q��x�Gf�5�AW@{�-��LX�d��փ��Z�$�|�t��u�z(t�]7C�ua�Q�t��>l̘�9qaD���5:Ee��LsQ����.*�xQ�tYr�$:�!yAY�������H�#<�]��kK��&yR�ч�,"������Y����7b�J��i�#�m�zEGN��u[9��(�C���)����ߙ.�.|j>K�:Q.:K_T�|��m%JoSī�Vb�<9�/�g� '�)��±/��~$�������y��Cަ4$*�#��䅒z��" �8�O�c`ru��$��2�+v�S.��gx	&b�U1�=�R�{�\@��:H�'�'|��>)�"��K��L��������Zf:=�!B�0S
�.(���VA5�KG�.����/K�~:���F��rx��R�q��8���k��<i���vV7�Zz�?-0(�1�Ϳ�#A�ӇM��+�1���wb&�m�`r��0�U(�e±�^L&�C��F��T�j�]M�_��~1qQ��A�{��Cbv1X��k�0�!�ב<�S�5�I��A�R<�
B����?ř�5�����ZKk�5N�#{��05w|V��e�ZQ tp�٣8�)S�A��/��[��ηN�K��Y�=�&	!�r
���v�"�?���gS�`LWt���mȨ���r0��[Z-���! �Df�{���Q>[����[6K��{�T��B�A_q5TD�:�4�Ȭ?&���f,5D��:z(L���QP'<g�8ը�G�C�L_�� �h����|��9KQ��Q�u˽���S����K-V���T3д��BmTd�al��y���-FSwh��L��nSc�l��X��;Y{���B���z
}���C7�x��.y���&d�N1� ��]�8&�U1�|g왁7e$����s���ќ�7��&�7Mk�F����B�|��c����.�Qd�j��Z#:���F#�A]���w����ˆ��6-ɦ1VR �l�nk�r���w܉e�޲$��+���HPQg���n�����2����۪-L���C|:��i�cA�יy�=�x^�Dx�O���z�u����:m���=Y�f�+��q�-�j_�ك��/zMҙ��akMX��,8�q��%μҪٔ��g��M��OL�}��K��Ɵخ�S��\/��5��s�mDդz�U<�5�#��(J?^w�