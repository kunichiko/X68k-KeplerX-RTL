��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#x!�S�q�x)��t����a�� K,��)3J}���d0 t���NҊ��YkԅE��~hG�w�Mj��G���Nl�J�r䛷��������-k�P�E�3b�vh��偍>�Lc�T,�`�q�,����ێ3|�dQ
8���l�h;4���?	L(b�E�;����9��6���x,'�:d_uK���!<�x}��o�]���V@��0�jƤ�Z|v��G/�"2fڃ���J�Y����ʾW^�1�z��C�:CvVVx�cjw�!+��-������;��~�r���I�ّ�*�v�J�y�[a�9��ԡ~��d�7�Z�y"�(0�N��U��)��Y�HE�
����Yx ]�����fiN�8*L���&F�N?���2{��8!�A�Lk����}ܚ�ٽ>���r�`jjh�S/@�:�#���Nϋ�7(�?�{�k�g^���|nv���/!���� D���|��=mY�{��W��_E�=[�x�)2(�7m�Lwr�Ȩ��M3
���c�ӌ�=���FG#TS��H����)�7�e|:4�]�{��s` ��n.�G�i�D���,�]�澧qgSB�L���(�jd?0Bay.4��\�5����-˝x�&�����|��,ߝu��
��I�BT�?&�@U�I+��5����%�C�6��*Í��k�f��f�K��F��b�����cH��Љ`��LX)�-7�n����*�f5!�6��#�+]�*���p�c���(1�@�y�m4�j\���%��6�l�]1k��.�/NN�Q4����6(�@�jf�
(���=�փ!:�]}�ə�n��H����Q�Q�U�V��yډ�R�
\T6o�z��J۽#4�@�|��O��*l��y3� ��R��5�n=��ӂ|�fv�Z�&x�%w�0ڝ�>�`��-�.��}
>c��k���۠�"��3����7�l=�Zl�B�S�P�����+!'�M¢x���(�*U��\1e�o˜��+V�H��4�%�؇�a۲7��G]��G'|;s�iIq���Q��Z�ΑYxoW:ך:)z��3:1���V6��	���WԞ���W]m۳��Jf�@	4�=|�����w��9op�nQ۴���`� �悥���Ǎf9�qջz.O�2�O,�a�䒙��������݂Bz��"��0�_�w�]�T���x�"�ڸ�?��4*,�Д-ř��"F���.���Þ���|�Jπ�[�a�!���h�m�y�õ�f�/��0�)lo6kזWb�
\d��S��)�pgN�~X�6�T�
$�bl,����In"��B��M������9�S�S�E3lW��t|M$����~NO^5�D�ם�`cG"��_J�e��}��X"�D�):���v�L�@ς�ꃲDK��QeJ�+S֓��v�����cp/���R����w��ӥ|�a��Bz���Q��{l��{��>�9�ItA�,]F�DI����O�a����	`	;E<GM��2�u����}�>k����c��7y������ʲx�L���0��܆mI���-<Y1�A�z����+�][X7]t\�k�%�G�A'�N"A��b
aib��nUe!.�!Es (�-��������!��ʓ����ȕh�@߾ؓ�oL��f_0��	gLFG�]QlX(�u�¯�9hI�u��`��w��K�HL�P\5v���l3��A�>AZ\���E\|5T C�������W�dv�u��;�yz5#O��Ⱦ\]K�.�*����@��	2`��٣]1��<M?hm��-;fq"$]sQ��c�P��/s2��y�3�?�G��M��l�9F
Ï���Y��i�Չº돠�$���o��Ӂ���yY��҈,_���F�q��)��4�%?��p��3��ǱbB��X�Ӎ�+۲��pw���9�
�� ����MǷ��p���	}��xXCn�r�gQ��[�/�<+ˑ��'y FWpIƫڢ��p���3�ۖp��ʏkX5)��f<�2Z�r��� �9]���6l+�rd��0&Ұ!���2DsY5܅�f��dυȓ�x<fCw��(�O=��X��}�y�se��o_����$��Er6\�;���fs�o��|r�OE�Դ!d^��t�|jh��Lu�����Sy���5��*���=JT��h!�u�o��K((�U���$0f?$�k�����K����iN#h��۬H]w�s��m�C��9B�.��X�B���XH�#(���MQ�\5�4���	�3l�%�Hw.�+rP�ן1��}�~c�/NM�ޤ���W?l��0��B��e��|$үQb�,�g->��`�dw0do9�Ldg�L��n^uaA��#_��v?�u�Uh��-2���˜e<��Ǝi�^,�e���(uJk��5<��ft�*�r���t����+�B�L�~Ā��]���N� �$��(�-��y�p��L5#�Ʀc�	�Cs~�'�I��J7V��(�����M�e��t��C2���E�rAn�`�틮���A��E��ןP��(���]:���}�31�o7\���?fPt��;a����<{^;�l0���j��\�?[Ԣ�^�m/@{�P��9n �;���1�(��3�1��]��,?t�uwc�`E��1B�}@��r������NUe8�S�k�SAT��ԃ�_��4���3�ky,�ڟ/�@T	uj@u<I�j���1��{��_����ڕ�p��b����z#�A;�Z�>���Ъ�z��ygD(�NE���Y��*����4ZX��Ϣ�a�`<2��?��7�;g 4��JZ����� e��}��Pj�s;%�f�o4�����~l�����P����k�'�y8��<YX�� �  ��(,F^�˛��2�o�Q߅}D]�1ȵ*����1��N�S����<����;�����d�R w�%��oW�,�1p����K���T�lM�H�|�����vM �͐c� �qy��3~ߎo��3������C�|���I�I}d�ҵ-��GJ_ʫ�JދH��0'�*���m)6���bD6xX5�E3��vn�{zK2w�8�>|��RS��!����٘�8}gM�I| �5�Hw��1���͔/���7�˯�oR��_K�Y!(k��@�>�[�^:��#G�\��O�]�1S�~��Ѿ@,�BG���~|B���Z%�D��N6���@�=J��ʴ�ى��9J�zn����B�z/|.��5����kN�����_�C�+�bN��ۋA�B�a(*����1��*?e$���2%��(qm&�)���FF��rY����@-~QTGI���̗Zg�����t��P���(��7�V�$� ���5l���A�{��~0�ձ�!e�d�-ޒ�����n�hTtS�I8xJq����WY��'y o�����5ϊF���d�S�f��_���§��LKźVm���L���Z+%�=�|���v	�z�嶏����DJi��}
�0#��PC�w"�����.����^�8��o�;�6�am��N�^��K�f������xWg��@�`t�|ݵSF�x���I&�Н`�+n�#�7�����"(2�GH�=_l|H��ݚ�$��%�H��}�eaK�%G>oIb"m�|��~�uӮ��D�ߓ�e�S�E�R���ݚ;��xoF�bfq
;��#�t�v�Jom�)���=P]�٤FlH�=�l}����������4�/'�ʸ4�D��Ba���%ky�w��Q<�{���gI����
�{v��([��a���Zus�b�3^���V�mr�;+�7�E"2���k�tų��#߃dYc��V��������T.)ƃ�8�w��y�uF���<�l�:����ǅ��֏X\B�]��=֓.(��d�޲�l-z�G�s�ͽ�7���!%ĺ��qWַy�k��*}�.�7�N��hHT1 �5�P����Jk7ۤ:�w��@<?k�O�'-U:��P0���}��2[,�U9�	��p��q����	�́_��@ƅ�B��Ed(�a����G7B�/��;U��' r�h��Jl��y*�,�H�+j��6��詗���a;szt���[K<\��x�=�P�CO(���y5��;��<Q���8	���2��������yO3E3<���\�%%J���8Q0*J�jE����%��\:툷�T~��B���V��A��8��X�x�����Q�����P�f҆����b�ۄ�3���N��O