��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�Tں~�ImW�.�^�ᆹ��������]��%�wx����xeՍ�ϡ�&JLc7e��~�'[�b(�Z��M%기_��H�K%_N�kV�.���a�����F����B�u�E�[�D��*{2<(ڡ�Ki�x�$�u+.ﶓq{�S3i]C}��}���O?�C(�M��:�+i�"7dѫī�pGKW�nvD�ޞ��A���1����m���ra �;'.L���c���JXcr`�����r>�LzJ���ԥ���H�q��ʻۙ'-� i�X`4�cck'g� ��nU.���!dj��(��%�\k?؝�-�q
.�X�����1W�`M��Q?gB��@e���=�����`ޒ���B� ��b���8��5t�V�w�`/4R���ĵt��Z0չgH��[���b���d�4�%�.W�i/湍`o(Ј[�T�2Bn�O�	�����no}NH���+�OE���]��ֆ�@��>���H�P)ok�Uz�s@Mpؑx�{��RQ��P��Z+���C��1(ꠝğ���P�[f���/����Z�-��?剗'>������c���ft��<K��^�����9G���&~���(ĶA��A�����<9$��ٺQq��74�y��jaX�#=��J�A7�=���BE��|�l��,�C�'��A�����)���S��O�8|'�6�eb>k�Y��F>Vs˼��_���X��p0$[P�>�D�t��-K��Z�!���=�T�Ƶ���+�����n�I/*.�}�$\�6���̋��!<��:6�Я�g.)�@��G"�߁���
���X�ϞNr�~���8�!�D�4P�Nq�u'��6�g���\y�yv�.��2�~���?_/�:B��Pb7gQx4<'=��Q�Q�e{�������D����Q��F!�o��ͣ�[+'��(,���c�^.��H�ۤ`q�q$=(�R��F�v����s��/γ������byA�S�Ч {3M�B7׽�܆Q��P�a$u�8V[y�b�����c@�cN�� ���;>j�r�H@�񰱈e�˧���3V��5�!�6��٠�k����%���k�9s��}���>پ\��.XVh��k����Y<��a�7>��,�k���l��M�Ƀ?
���'!��,�R����e_���KM_Y�w=`k��n�"���S�᠎H��Y�7�m�����#��P���nQ*���	� ��!Y��)�T�S$��^P�ٮZ�Y4�c�/�����9��?p���Ci7�/1Da���M��u&�j��v�|�$O/����6�K=�3>~���g�d>ݘd���PI/p�Qރ�i�	�-V��[W\��n[���t*(9�v���5�/%St:#��Z4�.��@�Wo�}��AW�N���_����3��h�xe���}U�n$�5B����_Ӗ��5��Upd3bL9��x�j}�̊Du[�S-��Q��W��Q^gN���g�E�����?�=�2�F���ڠ��+�M�Xǚ���z��~�zTj,�F�OD. <ۢ�]�]<�� �K��������:�����N~:>��
x����H���h�;/�t�A�v�)ژ�)VP��Wkw����yy���ި]C�����u�F��pG0l�j஛�^>�6�����K�\̍�����#+i���7yhK��T��6�Z'���m�V1U�V�w�����j1f��� ڵ'�]W�Z7�����,��E� M�K�:?о��� }��&_e����~�m�7��=�v���R��?��'R8T����1)L���8�B�$,���D`�b�$K�G�2�/ײ��`��r����,1�L7�0+�@��G/��	��q����K��,��������Ƭt�!S�g=���$i���1�Nݱ�/e�p���Djv�ZwsW�+��+�Q9��	j�2���!rHbV�Eذ�-fn�
B�H�0��g���F
�*5Z{G����Ƣ=��7����'���
���::b����ٵo�Pz���ϦG�an-(����P!��?�}8��N��m6R�)"��D���}5o4�W*R�VB���}��"�{*8�w��-rP��v�"�5z(J��s�t�7��)�~����:����,aqe������b�,h�uI��0K���20?> T-g�\s���c�(4l�*����v���_go�ǣ/�d{vg�/+�a�o|�C��2��B'����|D�g��ׄ&�V6}5 �2,j�S�3�N�UZ-"/�����N�2k��|B.Ŭ?�/|rKb�j�3ʆԪ�?E0lk�"ZwHB�g��'6����U"3��fb�LG���MI�����F����ߢ�x�����K)�Y�7 �xj$)|�H67�I�%eɫJ͈m�C� ڤz�{\���ykX��i�S�E5�x]�WN�=3��A��i���	�eO�cx�8Ӓ����f����d�']�]����WМ&�,t�%n���N�1�����ܰ)�b����{�O�����g޾A��
Ư$�y��rt��5�]�h&#p�ni�kj�=�������auE��*k���a��&�0��a����xzW�L��ו�k��s��,��Ӛs��o���zr2a�fo����I=r������jc��)�Ym��@G�.�*���r�L��23k��{3�x��;��?߇wڇ�3����8�u'�4�l0�rVM��ddB!3D��9�/�=�1�7�c4C���f[�zO��ɉ��4U�\Vi��t�ϑ/a P�|�.�g���BqЬe�`UМp1�N{�5���y\�����8p4�0�\̛���/{Ē�q*"�.R�Vx�%�8&C#k�ZK�1�O�g@�ŗ`��t��Ln��3t �^����9�E�C��� a�,z)h�ٳ.��D/8A�4�	�l��Q�p��g���X���)J�txFo1^��Y[�E����Qފ�\�+��@#���EL�;�*X1��-���7��x�E�"���鉪V�8�4��׳����ۥ�ҷv��t���,n&B���c�e��%�t�d궣�ҭC�}"

`}:�&F����gt�����LR���cʮ��{_��0��Ρ����W���n��X�!u��!3�0��i���⩞��� _�l,9H�ԙ>[g������_Z�^~����S@HX>h�p��X�I06��iL�b-]�����
�>3Hլ#E�<�+�.�"-�:J,ِFj��9���p�/�O{�>9��;�_}�E��0�7���7H�dS���:^ؚ�e�a��+5�0Ȼ���7��W ��Dǻ���:o�2���-�N&�����l��6�nv����W�m�[��3�z���wǘ�Y!^���N| ��?��!au�xDW;p��%?1�	�>9�EJ�,
2��wt��|d�ZѴ���べ	n���-D����N���fTmZ�mN2m?�Ph�c N��_�3�COM�4�hu��NPP�(�����S=1�<��ْ�����jX��� 9��o'�z^M;=/ ���	aSA*�h����Cܰ�@8]���{M�dX��<�˴�ѓ�}��f��N�^-�z�ug���xE�����o5-b(�'5-���H=祖��Aە�}'�0���_D�R*��SkW*߃Q
����6��_t_3:��x��	ytMB��l]��6�!�|�M�����v���GC���(�}��H;��:/�X�����v��{����}���	��4�jŞ��
�1E�Dt�?P�H�҇�`ɫ�\`݆m�X��}��$��
��I�rX�S9l+q�>�V�̳�C9������f@iAV�@ˀB��<U�V�����,g
�*:yO-b*J�cV|��X^�rW����@C��f����ڔ#�E��D<�V��r�=ؠYa?|���č�>�]o��3��)��b��O�\T�l_��ZF�X��G3����6����B�|��!�ABT�"8��w�~���Y.���U0�=z��X�F� �-��$hS|>�t�
�)����	]*��m �c�/�[Xy~Q��:"���-��w��*{>�Y��C��u��a7/kB��^�1�/хd�a��_u'ݣN̛��kw��Y1G~k=����0�k�r�K&�-�^_��!���X3�"��A�`�z��T�D�|�I|�IٲfA/ڭH
�zH�>`��c!���ۗ�;�JE?h�յ�S戥k�6E���'"�ꆮ�����j<��Q��m��o[��l�E�����dc(4N]B\����q����Ġ���QyyG�#{��[�I�����)9��aE%E"y֐5T��aϩ�B���bֻ��=/ꮄ�0AJ�y�T�5-1�Z�A�� �kn��h�$���T���
Lh���΅/����#pC'b���δ5D<�%��J��@��N���#�Y�\c�z
�G�O.����7��(�н��93��d����VP��c���+�gF�<�@�� �A»L]��O@���"�<���c��]�kYv��$��1���� �2�x%�p�R�E2�E�	��9M��/_�	9:؇>�F�)�ͮ-�v�^��1c�0e�w�j�yG��eW I`��?DG���g��F���G� �):GLt�U�ץ>���DkXZ�109�*���r���>��-9&����A�T�7��w
��%=y�
�4=ѷR}�_�~CC9b0�.6{&� bK��K^5���l��� P��nxJ�b^���8���r��	�m$�A��׉̕��Omey&�H��'���<LŏJ��k��م�����V
$z�+�X)�'�������s�{a��Rj���[h��BOb�&	�q{�,�]�[N�J3��tr�>HNE��1����-*�E�rWN��_���ZYU�]La�H[L����=��MA�QJ�A 5��z�9as��6��&vq5�?��M\o��d�Ma� ���_t�Z����Z{���N��̣���;Tp9�̄��Bgn֡Y�CY��ۯ�mx�#�Yk��:�C��=F:�9��d���Aas�R��V����h���@8p�eN	��S/�P�M�>���1 
`�c�伲Dfse�!B�s}0���q�˿ J�Ji�D0�GL��+tJ�D��!���~Hh�Ř:W�`ʋv��x?�ľZ����,��_�T�ॳQ-ɲ=�]#�m�)WEY��5�by2G�O|���v�?�D�q;��ܿ�#�����8ڰ6��!}JUIG��֔�ř�M�I#w��VAP���.Hw��:E�%��4P�gP@ E��U�1��2N�����K��������1�!,K�(wJJ�Օ|b�K�2���d�,�*����`C�e���0�(���C���7Jv��-@��ߘ��I�{Z��3�P��7p�0QK�-&�����Ӆ�{�.���	�%�`�3+�4�z'�}ՃÄ��8 k"�ZC-Y՜v����_W��ߘ�#S�Q!k���U�nh����<�7�n3��FD�H=�)�j�'�]�ӤýZ15l_��F�����7i�7�a{�
�I{�
zZ%V��Fvj������>��R���9�����7����d���sИE`m;�=��ݸ�U|M���ﶬ��V���r�+/
jk�;�G3(mqP"��X��I�#>q}�tuN�g���F��)8�'eO���R��ޜB��b0&�3��(�'ec��|s���%¥^a=��L�vY��
��B��7�}�J8n���4�ޣ���q�z�����������L���(�����״�&�ܵ��9P{�B��@w����n�'=о�E��O�0n��;����2Sc' �V���#hk)J�'��,�%X��䆹>oq�++2]��z�l�Q���]��Q�䠝1������*���B]m5�X~)� D�)��? �\����h^�:��2@���"�q�[����̧Y��U��w�X�ǄY�-NX7���x�<D����^"z2�?�RpQ�3Ѫ�kx���_�i+�i��1"B�9�8�Dg�jcO ���T�)����>B<�!`8�QN	B��l�]�k�?�e���Q!<���f�$@��=A���%��e���G���|�̡%��x��v�[;$`�˂U^k�o60��8�gjckt#�����ATH�DsҚ��-z����r�����*����߸
�	�0n8Ժ�ǘTf�رl~Gξ��e=��y}_����4���Bâ(��+�88*�;�k.��ԧZ�"�Y.n��4��(nr�ס,hV&�f,O�}]�WmE����wYZsj�<1�r*P�o���2���S�Z.-����TD&�^���`�-�8�7�nh4�x���j������}岰���"H-����h�E mc��
G�m����n�EK�����9MX�D�����q#� 3�ճ|�f�w��;h�e�B�]�E?[��u�2��%��3Ӗ�s��쪈���<�L�����JzG�f�$%W#��*4Ǌ�}q�(j����NEw���m���m��^jQx�P�c1 bA�̐ ��(�DH|tᬍ��Eݲ�إ�9]e,rF� �H�odMI���&M6�e�\�\h��b���
��`���F�_`+)��M�c�ЕSح�O��rV��n=_{���HF 6nճ@(& -�=���^�ĳ�+����-�CM��H.�f��2���:� zS~K��s����ε�{5�y�2~�2��_