��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D����gP�������������44��Pg��w�k�n�L�t�=�ʠ̲J�=�	�$tG�讧��p,��sC��Xu�_ S�	��mZK�qnu�*u"ǋ<�L*�2S���!��i�އh���
������)�=k��l��hx��I��} ���l��CaoK^G����F�HE���}�-���8���C��)�6v��q+���BɃ״��0�Ўl���Ax�`93Di�j�]��0x��uHo8ȁ�h�+���]�,L��uS��|�>5��9�8>�U̒ �|�o=���{�
'�[	��ԄgI.��Rs���Z�GݲB�_/h�_g�ˢGmYAa/E���,Ӥ`�΁b�d�@��+
��kz<ˤ(�w����0C݊��L87�C��������z��H�w��ڻJ�:>A��>I�B	�KW�-H��
 �ѶJ��;�\�16Ji�,�z}�:d�9E��_����Z���o-�[Ɯ��F$v�KG�%Z�:�oA4w�)[����:��z�X�o=B�e|�_2��ͰUSo����I#ظu��#x	oC}�v�%����KBU�2 p3 e�+�0ʝ��l�;$랉�A��t�h�?\�<��d"]���xuB�@3�{��e40/���GC��������ھΛ�HWR4��M�q��q��x�Gf�5�AW@{�-��LX�d��փ��Z�$�|�t��u�z(t�]7C�ua�Q�t��>l̘�9qaD���5:Ee��LsQ���荌'�^�� �̓�4��QɊ��������(G��7��1J�dy�>� ��ltOBU���qj}EB�N���紐Pe)#�P#�ٽa��Q�ܐd6l�u��=lIQ7o��>/Al�c
� �*�wh�n����6~�+9��Q�*���t�O�@��߾�gdD�g�e$ݔ����Q��d<D�n�IV1�/���Fߔ���s�L ��	��qp*� �x�k�@e�(ʜ(� ����jC���p.���1���LC�*H��U�,}��z~ݽ,����V� kkh��@yX�[��+e;B��tX�01���3ͯP)��mP�S��Q��������PЁ,��0��:T��y1��+x��r��������D������yJ�apbK�M=Db7BI
��n���X$��C`�����Mr�͔��f�n	�XM��2]��kj��K_@bо��q�����o ��$<aYV,����B�z:P:]�R޸9�?�Z�*�*�J}`f�T�-�c�OT����K	�߭�ts"ϟ�����w�=���=�̌����g)�]#?O�H/�0�b>?����h��U��~�c�b!ا���n�"�mA7�z�oI�w����]���k�ˬ9���/W��ny��Z�Bu���A���ǈ����׫���	l��3��h�o�g{��I��y8���jMUOsDa1�Yت]l��/�<W�&)�#�BXL6S�/X3���Yg+ct�%zP��7Ϟ���ٔ&\T���O�4
�5�tr���`�A��E��������ټ�����(�>�3#�X��G���5'�K۩z�',�%����ݮ�����9"�X8.���q���\���z]�bk�"! �����V+A��[�>�Y��-X+���LØ���R�G��'S{x��p��Dp^ݷ����I;��zCt( �!t��
�ni�=�Qh=�_%1ጞ�i�x
������X��T� ��r|�7� �2�:�Jw�M?�sg]Ssfa�'�;'��3m��6m��K<��]��o���B_[���٣Hи��R'`�J�H�$p]�]$�G��!���뱡T��-�+��i���}�Ƽj# �b��*%��?�~O��/�17�Zh�ld���TL��>��A�4��?U;�╍Hv)&���W��>(��a���x�ϿRM+����ft��K/A��Õ��*xw�2{<`��O�h$;�� ō�R״C�Wѫ_�Ci�^Ŀ�2�
@g��ȗ��q�"��`�^h-�:~�|�Mv�z�_דNsOU��W�s�������N�˯C`��{do�hLph�9;y�SƬ$�{�u|��+T<z�j�87o��[[��ŰP��?AD����4|�?���=�2�♡�bJD;�����~�(릁�R.���3Vl��h�Ɲ�����GyEd'�����U�%�	�$]�R�P�����뵶D�ݑ�q��h+�b�nŊsrUh�2���}\�Is�]=�z�U ��j:1��?yZ%���}�6����$��)(R2��sh)�S�O�27ģF��k�e�D2�|d_��#^3��̳��q�����>�If%�?2��Ƽ�� yc�*���������=�q��`4"��ī��4T:l�_{��K�w�F3F&Ļ �SO�>�{�I��Ӕ������h����6��ig��f�8�d�	��D��0�R�/R���c)��!�v3����?BQN�l�L�!��ŵr^h���Q��D����6�'���z,�ƢV�.��U.ژܡ�੉S���A��**� Z����u�8��D_�SUV�Ϊ9|����	�Sn7t�g?����Z��{E�H�n."�x1�eܯ����5�Q� ��z�Ǧ�,bʶ���,�#����N��J�Z~�>�C��9�VL֒����Q�|�]t3E��`���G�6��{D[D<�f���泳P�1y�Q���r��"�������y�Q$����^�0AT�w<��;�Ⱥ-���4ޛAK�@ys]��