��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D����gP�������������44��Pg��w�k�n�L�t�=�ʠ̲J�=�	�$tG�讧��p,��sC��Xu�_ S�	��mZK�qnu�*u"ǋ<�L*�2S���!��i�އh���
������)�=k��l��hx��I��} ���l��CaoK^G����F�HE���}�-���8���C��)�6v��q+���BɃ״��0�Ўl���Ax�`93Di�j�]��0x��uHo8ȁ�h�+���]�,L��uS��|�>5��9�8>�U̒ �|�o=���{�
'�[	��ԄgI.��Rs���Z�GݲB�_/h�_g�ˢGmYAa/E���,Ӥ`�΁b�d�@��+
��kz<ˤ(�w����0C݊��L87�C��������z��H�w��ڻJ�:>A��>I�B	�KW�-H��
 �ѶJ��;�\�16Ji�,�z}�:d�9E��_����Z���o-�[Ɯ��F$v�KG�%Z�:�oA4w�)[����:��z�X�o=B�e|�_2��ͰUSo����I#ظu��#x	oC}�v�%����KBU�2 p3 e�+�0ʝ��l�;$랉�A��t�h�?\�<��d"]���xuB�@3�{��e40/���GC��������ھΛ�HWR4��M�q��q��x�Gf�5�AW@{�-��LX�d��փ��Z�$�|�t��u�z(t�]7C�ua�Q�t��>l̘�9qaD���5:Ee��LsQ�����yEE����7��W�E���p��~(��ZI�Mm�RP7��(����~6&3~ܔ^�-��=��[?���|��Az�_�^?�/�Yķ��������k�#͢�t�XW�@�t����?>B�L�_`;I� �Z"��9�V���� �����~ưu��+�8ľ ����;���$Ee�OKX@l�o���c7����O��R��X���:��m��6$�G+�4���-��<���)o!iT0���������1���h~���'�}����P�_z�gMd��cO&�*P+H.&�/k�~<�&խ��ՍC>��������/"�Ǜ��gǞ�'�-cZ�юa�s������y�9[��9y!r3�O��EU�v)�e~^�W��Q��=��H��ֻu��?.��NL������dF����`�����pVNuQ\�9�K��d���Z��rυ6ScO���r����;�.��j���a���3a̢�[e�xm���%��f�L��p������c��?c6Ӭy%������l�[.��%��]74][F�ђ/� p��)�G��P������q�_�:�"��'�5��1�Ye7pB��
�E~�:Yl6ΎM�T+����+y`�}��%a�qi������k"����O;��y&A&	)h]�����j�?� u���]M�ُE8Ô��t������xDq��0%�ËX� �5�E�ĴHFa��������� 0.Q������Iʚ��{pE��k|R�U�)�(�gS��Ё�D����Xfq�<��#��Ј��Ӏ��l�Z5�[9�����E����]]�復��h��}6��ڳ���(�aIbJ'^#|�@wEԡ7��v���s�v����x�d�����0'��
bvP��+�zi�s�~������⁯4`�t�,����f:�\+ ����x�h�Cq9�?c�o��q+lG3��~D�F색&���m$gw�[Ϳ�u�Ȉ#��7L�md~��|m��L|����x�E�'��,It��S��_䆔.	�	k-�ȍ�f}O����"�L5�p{V*�+�͛����h/W4��D�c�We�5>����VEl�\�_�cyt�;+��Y�Z��w�:���_)��#ۺe�+�����Z�q�� �	2#��e�uK�v뛁�5� �w�i�����Bő�x	ܐyO��j�J�d��r������&�9XWKT�~[���۾��8�eH,��v�='1{�yO�oDY�U�3�= �^��# �䜾��))ә���`x�N`������?�h=	��I��:Ηr ��)��β{��L����-�z3z������{Ƚ�:a�74�x�Og0��#\.g�_	��P���s���e�Tdl���(�ӿx��QU���˪V�v�t�"fZ �J�:X3y�Oa;Vɸ�ֆ�쬫q䁳~ɹsT���30���B$1}(n�v&��M�M ����F�e,�h谠z&>Q�
�n)�t���-���s��I��ɪ�_�� �A�xG��;]Jc�o����Ob�䞙��R:��Mf�mO)����F>6���nn��x�'�{P��a�JW,,�LyZ���+e�B��V���"6!�R�NF�x*�(����.�9��Ej�/^d�M�����t��ƾH�N��.���,F��0���D6��(�X���h�跨��	i�)�1>�Ї���f L��w�������@9�#��q�$���Uާ��l�s��voO逗6��n@�H���t�&�v�/VL�qt�ʳ�M�>��5I�57z=�e"�����hل�x�~o�[��6���9��,��'���2w+�~��ۇ�54O:�7L�Zz��*ù�g����H^->᧡-��~L�7�����"!�ӎ�mYҊ���P��C��kYS��|O����V�E�g���� �oC�4��K�&���퀱������*-b�n?n�DrRa;��*�@���\���V���]�ǉ-�7��p�"�
����㾄	E�e��m%�RW��������E��t~��̝���~
��U�Y���\Q����������9�F��	&v�������A��CS����2�&s$]m���@�F��i1I_���O��uyi�#kFN��-}�(�:����'����)�4��$�Df����k���1UN*�h>�}�[��o����W��	�5�9�qG�4Jl��1�>h�/p�|���i��mz��ow�hO9�v$T�&���.K�.|�Ըڬ���r���UR�05�}�ޒWm�RDe�X4MY�h;��ߠ�ܜ�45��=�/ʚ=�<4�D� P��I,i�����߀��ҹ\]�U2˭_ӆ��|�W=A��B���..��p�4�5�b1��ef��D)����*2>��,}��y���|x5�FT�e׼�U���*<D.E�r���ח���0F���|��7p��q�Yw7�խ�Ӓ��7�j(��֠�@�XiDvi���\vR^�ˤ9`�� }|��[�в�eR>����Gü�u�6zU�a�������28KF[�� ➉zVzЎm{�2�~h�&��H���}��4`3zƸ�@`",올}I�Xv�!�,�Dd|�����Lݛڌ7���ڻ2����l&��q�S�r��F����^��L��ͽQ֣�|2Ib���D~��[����:�f็�S��?���u7���4a2{K��]'��w��F
f]�i���U��i�o˜�K��C���y��.u3��À,Ƹ=qF^Ӑ�Q�t�c�Ѭ��IՌ�qF$���_��<j
Ή^3u����V]_�����^������_�Z�Ak	�	N;k,�>V��D%7�����d&5�����N���8�Z��{r���2�n�E��T�~����sA8���I �2����j�&�Y��l����6�f�7/-0�	H�3�����������"s�b���e����<T�;1��`�����Ɔ�4���q�S�IT�K�t�Gc�<��s�a���-�M�ztUɺl�1�S��J[N�A{f9��W�v������5�rF�K5GGE����u�5����P�8�cH���2R��j?a2,�齼t�̴���\]NR3�����*�!����N8��]]:��ۢ�X�^�)le�Ρaj�x���c��!Yo���蹥�A諞F�V�������A�s7$�y2k�6Coz�5�e0%���9t��3�"���y_��]�D~����Q��)U�}��&�}�/���4��	^���\���k��Ma�R��>ĝ�隷�J�BY���hoX��	�t��_�Pbh��K�D��o����uC��3���)NM8)�k�.�{?��J�Q�3�
�q�R���L�]5��]N���g^�~��tn��W���/)$c�X��a?�1RR���R����H*Ƿ���N����F�������>n:�+꠿3����ѕ���r�U;��aY�X�!�����٧�nk%�+�2���=���󺭇k�/��m�@��N�c��G�:��E
�Z��h's['h݂.��6p����p)�`X��˕������`9�v��җк���ÚkkL���c�U�F��;�٢��r��#�����Av��ژ��P��~1���y�
�:����d�u��
U����I��h&>�����j���!$o��ЕF��rΙ�j�8qa��%��4\���l�K [�{+�"���9�տ�u���#%�W�jD�E��=q��Ij4[�<�g�-p>tI�}	����z�f3Y��|�%0��.�+"�+�'����r�eF4a��Ir]Y4!3�#ފ���y��ۦ���r��=y~XC��tiq��[Ap�כ9��[�e�C嗧�-	S�|�&,wǡ=�����d*��803�%�>�@��YO>.o�9��G�p�C�6��-�pan���&��^ڰP�J��HX�����އ7�	�gs4f�����M�4�/7�����#7LGU��):��nJnJ|D�#�Q�?ggC/BAfÖ��
��:u���]��^<�c.WY:���:|m��S9)���<��B?��V�(���g�W,4@)c��B ߱N���z�˫���b�FD���O�@U�O� 8�r�հ`��Wff@���H�XJp����:����<�.Q ��v���B��wM��Q^�|)������^��˭�ܠYYr�gV�՞V�B������|�Y����Ŭ��0���巪㠴ߟ��*D�o���f5T (6�J^xf��נ��%s�����a�
��z5�v�c�h<
��E���椀?��(�6���/����Z_�*�_���,C��I�q8�����d�b)�|�.��{IY(s�������*�ĝ�=����efP힔0OV���zb{����fܕ-l^�;5�L���d	��M2����Kc�A�W\�&����/ ����G��#d��ǔǍ�w�5�B�r�?��XR�(_���+�,6�!�-7����W4��"��粎:	��ej�	D�x�3�5/K4'��4���!2�������ש�_�=7Sv���:}���� e�KT-e�5�޼3����_�MB�e��*+�L��Ƭ�pY)�P��2��"4����u#D��R)��!1��|n�-gc"?7����%��%���@�;��}����qb֋_�])�.%������# LiQHX�M������3��Fj����I۝ .W~(���AW����+nї�>Ώ�o��u2�TVV�ω���+���';N{��8�d�3���h鹟�ض��p4}:��������F&ƌ�a�)�w^����;�����m��ػ��V�`��W�!y�;.Fk�g紒-+������HW"�01�]{�U&��깖Q�˦�+���	p�#�s��؁�>0���Whg�ZT��#H*c_������s��"ѰN�`�^h��Gw=C����������s����tM:|��C7i�n��r0���=Z �	�����[/����TF���s%�7�V�&���,V�/�c��Hynr?�ÙI�Gu�؄���z�S��R�3��{��:��))lߕ���8���k[Jͫ�X����Q9�Na@o��,�E�`�'l�,��.��A�d{�b=�_e��O�ܑ�W����dKm�gg�K�N6vD0S O8ȡV�_���J�I��l���ԨQjiy�\�K7,��P$%,�!ǅ��P����B鲉,����7�
����(A}�ޛ���
��,�����W4����$Gj(�\�ps�T�4��=�5?�6�'�RtT�#
��y��6}Tm���eΞ�/G��<�ɀ���h��u��e�*����z����p���4=��DP��9�q��g�$�%��QqG\�.f���g�(hѧ���A��4�[4����&��G��ij���7ZW�_-��͟	���U���K�3�}P�ޞzh��7�^r���Z��	�.�@`G�{��Ǝt鿗dr`�� �ȶ�O�/����[���* ^Lېe�d:�uN����^�RR��3�ڭ붊�N�
W�����W�e��92=K����M��!�đ1l�K�~u�4��¡���&����cM$3�B ����4tр#9�P�tu�^���x?1�>5�2���m�������a����!W��R���,���o������U���P�ZDb��I
��$+@O�(������ݹΏ���{��)����S)�x2��Ё5�}5�A����ťVi������J:��%���߬w��u����ۺ��T�����F�ң�&��dQ�5< -z]�Q�����7gb��`.K���%!z���/�b�ڋ�0��M9���p���V�kc����F&�m�(��B��b���֣�#�A`Bh���'�9�N�6"�,���v~)�Gg��"�w7��yu�n�M]3	�o
c����W�FDxP���Y$�+�D�Do��H��+���#�:H�6�9<�xH�� G�ȹ���ѷ}��r���s4N �)v��;��-�D���̦�|,n��Dq�P�Z3�#M8�������D���lGeE�;�h��qh5�G���[����j#^o?�m�o3�E��es������/�f���D�܋Q�ccN�&&�w���
�7���|���8^p7:�{�jP+�9l��[LSH�� �ƀ@�	�j'5��T����w�5!l&�lrz�S��f��#QQ�:����
b�ə�%�q�R��n�`���^yh��¢_��a�UV��x�p�^p{�����-l�Gj�9�O��q��c�"=K�8^�\�t�ً�s�G��@t�^:�n�0���Z������Y��9���8|���rZ�ϯش���LvOGK �Wm���}��\�;�yN�O	� ����<��K�ܬ�����ʴ1 7��(<��ӛ�GƣE��펤�����.�l-|>�?��J��r6�C�n�M&�GX�Js*Pҡ�-Z�����:���;���!_�+�x�����N|�y2��ł���%k��z��[�9ϲὦ|k���V���)�5���i�X�I�e�/�	g��ǖn[P�1���<�����TrHl�%c��F�}��j�������L%"� �-��h��믷��VC�����)h�1)� �ѕ|w�*T�wƥ\�ֺ�ӫ�.kC��}J�=��qI:
{b"`�ޙB�H����q��G�v�;�%=Z������R?<�<xϧ�=ol�ӿx����x~�b} �u,��e��
}K*B֘�@��}9�/s�tv%�U�M&� �,��ܚ%[�pEmC}s:�d"!Pq���>�����̾����_^�h;f�"|��V���)�^5��4�'�UC���5�/Aj���(��e)�����٣�r'��}6ȨM.���Ӝ���=���/�/3qv�b�z�k������
�<%-W��K�b��
�C�<��\�s�w�%E�E�W7;/d�has#j$�q\�B5�VR�ϩ����_�O��ȴ��$�9�c@wꌔS����1���%l�;4o��Kuχ�V6�a9����npʢZ��v���y!-����4k��>2A�����1�\�9�q3��%a�b좥4;�. LE5L�
�;���vnAyav�o ���� ���ݍ.�a�,g6Y�R赻�tP�o3��lo�����l4
G�BƤ�O�Z�F}#�|^�f�/�G�n�^�k��i!��F���[�}7�4��1P$�Y<e���K�@^�\c��+MR�bS�h�:��q�;�m�e�LƄ-��xjWNa.÷Z�2*3X�q�k|$"��@/�Vqq�&��7@>�<'����3|O)����b��N΍�7�f�Y��Q](�G��T��	͓o�s����@<�k����6��.���tt�w�{��o`��J�WAŏU13}O��Z^��V��Btm���ﲷM+n�v������\�ζ�E��p�~>ty�|a3���p�v,� B�q����]&�sW�J!ō�\U"/�^h]�b���=2X�WG��@���q�'�U��t�x�V��9�e�Rk�>٦�xy���D'(���%�����[���t3�UUM�Uǣ�z{U'�]*����(���&_�ķ%0Bq��@V��CC����%#�p���ڠD}60� B+bI�QSX;Hm.J����PLF��kP�'%�up��̹�ha/��Ec;{�z^o��bz@TXZ�pP���
�^:l�Ys�'Ĕ��0;E4�]㠖�S}�A��%s%�A����>��ȧ�vTt�l�|/$�8�1k����	��9+�����l��sz�n �	Cj���1����pzH�uNN-V.|�#���v����Az��J������c.�f8�^��%����c�/p�C/c'��V�h��{�#M�����.����̬��*Ț�b��dң��Ici=�k}D�囍f�<�&	c闁l�۫���7J�w�j�iB�Iy�~ѹ��R���i6p�q9��n�����.�t���B�Y�aA_"Q��X��V{>Ԑ�cժ��$�Ϳ����(?	�-1A�^�q<EA��[��ҏ��zmć�)�j������RE����6�M4Țto���U�-�<�'��-�"� �YOꎣp��F���HQW�g~��˗󏨞L���$r ^����	��p��7�������Vk��a���d���"f���?����=��1 ����y�Sp�~t�%���F�Fx"3]�����ut���I=�읐�Ka(G�ȱ�t|�6��'��<�r|�Si�\�@dXK�ҟ�$�o�����M�P�G�x���]��B�{�M��n��h�Hg�9ڑm�ڿ�J�'��ʒ��y��W5)���}�"����-����,�6Sa���o�)F<]�����TI\�pD'���q$�M��_O� �ą$�l0r��e��i���)d�g��l�Șr5߁\͇�[m�B��4������3Q%N<�;�i�����-d�CN��ш� 1�	Y���pk��xj-.��&J���(��p#y��X���Q��-t+v�H��)�����@�6f"1l/���3��r7i�^�N� F4ޮcؓ��,Y�۷_+Gfo�9��T�ի��qQ��D��+?w�-1��F����P	�я�ڷ(�%v�f�o��W��g�I�OV�*�M��</�=�Ẹ��!7K�����J:G���"d��hdc�nm|���V @a��KG`\5��]�Y�n'9�H�0�!��у� �=@X^�.���`^ތS-9��H������n���h�q��\��w�6�W�?G[
r}|�ߔ�
������,�`�f�:����o<�����ƷC�-vۂ����n�|��͞R6��W��]�M����_�Zv�����*B�Y�V(���E O��d��x��;B�!�Mb�(�;�fVo���(v�Px:����.kB8��:�����TR8��n�L��� ŉ���5y����ƨ�� RC]�&=�����O���02HE���)���(~�*q��������-���1�n:��ecZ�I��1b3j��&^l�%4�X(0&R�WoߧPpJ��W\
�'�'t�sqPO�i�tM񝳻�g�*t��9�'��:q5?��c�q�����CZIN���c� �]l��YgY����s�n��>,~GK��c��N4Ҧ��Rxu�{7�Ɯ�{Q&���O����D}�v6�dih�
W,h�E_9��wK��K�W�>��@��@�jU����%�mT���8��ɲiq;D���.a�<����6� ]{�5��αϚ��2��-��}-q�)ղ�nj>P�)�8��̊0��0+����?�Q���y�*S��[�uK�y�C�Ŀ�B�Ī�9l���6�ix��a�VN"����~n��1斊�{ҋ\
w"�f��@V��1l[E��VT�o��rv����{fJί�f�����fȚ} Mz?�"�E���c��Z׻�9jI7S#m�����(�o���CD��k�,a���#�}lL��k �������(1�=�2f%��� ���<����sdUx�~��G��6�����,���g�l
��n�"s!a.P�ߐۯު�t�V�*4��>�K�����-�0N�o���	?���)H�H�.�ym'�_S�5v����f�����g�	ѭ�}T��y~0m�z����r�����P�V7m26+���L����\|O�6k��:����$gǕ�Ǖ/W8�̤6=�2m 5�����H->�aeH��6 PF�ھ1�r��`�l��=RD�ޫ�xw�;5����.�N��G�n�5qI٥�a�41�6����U�_�i8��£�>lͦn1޽A�`+����P4�m��a;+S��G���V�-X��mH��'���4��%P9�Zx_`�&��=�V�	�{d2r�Ž�2E���t�\��Z9�n��)NTE@��<��s�[��dr�Օ�ʴ�6�m���݇�_s�I�3�l��~��W'�v�`/\Z5e�7+���}o�V�4�Uղu���F��:���^���"���7����8���&R��#�@�0�$����Y��[/<i��������8w�C��&�`($��f�B���8����L7GF(&������`@kם��`��nT�:pg+ �F�Iޭ�鑈��ȆA����lxۮ)�=W9���|f�i�����0M��б~���=��N��-�2��_2��H�r^:�@�єb��4Q�sV�4f�(�M`�;���#�%~}(��d�l\���T��rTi�ߐ療Y8Vo��	��_\s�1�����+T�Zr�ة�k�\,��P���;���\IEΰE_�B��o�d�X��	���j����p�w���� m9_�a�&����S%�1�b��-�=!6vh\��N�'��s$]�F9K�啯��W���dߵN�E�I��j`4_�Sya�����D���У���bf��_�\�����%p�p-&�u	䶤��� ��GH$��{N�5�8�1ñ�;�@��ڀ��m�r+��*ÇW���no��v�[.^��ފ4�^���U�����|q�͌�m�|J����b��Vp\V�5�*aq����Q�P�˧�,���3]��]�������ef7Ԅ��H�!G&"^���9>nɡz7ʋj�~{@w��x��?�C4Ks[2��J���ߢ�����LB�Ntϭ�s����-���G�6p�.�e�pql�}�u�`�B��������T÷�3Xo��p�?���C%�#Dj����� j1`�k�q�X�~o����>,��%�:�j�w�W��Ci�6��$��:�骥}���dG���=�C���Y�I��ZG�L��c��M������\��3_։��s�/�ُ��g�M3W��e�q4]�Y���^IdHs�f�<� :+\U���4�4�� ��|���}��1�&iL�݀]�P�b#�߄��힟X����O�8��8u/���>�<T�N�(�" ,�"8��KS{����X���p�$B�0�{����͂�����o��6��*�3���̍�M'N�9ω�0��35�(�7Jd�C��3���ױ�Fsa���{�uמ���$T�/�NK�y���N B����B+�
�������W����H���w����x���e�Zv(N��/�(p�_ű�۩\Ƶ�������6�z�5�*�0~����Ĝ����D~%1���3
��%=����6n݅��9}vʹ����uA�~������`��4?!O\!���&����fTr;��P-��F:��D�@ӑ��,���{�����1�Jc	�|�%�f,�0��ʝY�իd�>9�g�א�I�7 �@Lh�Eپ�	G:���z�7�7gʔ���#fЉΠc���ȕN{)�%�3۷ԩUVL*�di e�-֫h�q��u�a�l�(tF�ql��Ē�+��%��H3��< .i86�����p��ߊo�J���D��`l1ad{�L7럾�7p���<�n#�~�3�P]Y7�m�#��wI|*��>'ʳz��7��}�}"�Ϸ�<��+���#��4���lû�kPd�H.�ǎ�o�u	��8�B���8p?U��ZÐEaס��v
������\3��ӝR\g�~�W�
y�H���IN�,f_M��>�-n��\��	LA�"(��p�1���1�s߱��6��U���u��<�%{_�ԥ��-����U�̴(:��N����ѹ�e���,A�Rn�e����^8�|�f�� I������&io��r��kUo�ً�W�{n
����"K!�>ԒV��~z��� 0h89��^�?�A��z� p��~��a�DPm;�������Z%N\����ɣU͕2��GN��DMP��2EV��&4!.�Ҏ0eހ0R���w�hӟ�8������e˓�ܱ'䈎�&_
��Y�[�#GՊ8�dR^���2��h0�ڷ� U��=�{�.^�1jF��H��kk5��J�d�4$E1N~j?^C�ձ���w ӡ��Wg}� ^m�P�o.���
O���M�j��z�<�C���y���y�][��lN�/�js�����!d$�?3uT�s�~Y\C���T�&�fhh�њ8�Z9�+��r���i���wr�6������s+��l��O�!fc�кN!���'�>�x�H��v�0`�#��d��Dq�҉�|>@���V{�M� �Z3W���b[�x�6BO5U�2���K[{֖:�Y�S���^|3ɸ�^ �CYa4��[��X�z��qf@�>�rc��7)}+ �����y	�+�]�ߊz�����*�!vFt&�_�
�BD��Zp%8�%ڷ{�j���HKy��7=F�i����^��'#�z�	K�W�����r ���4�C�滑�8�e�-��/���%V����G3TaU�����A�ш�e,�t�Or��M��Z���a��(br�r�N˹�s,���q֡�����C����"���K��p���»�$�B��@�#��]�*�Jᔫ
����p�c�W�#D�ʬs=qB��<q���m�?��f׈f���q�f
�Y��S6��Ѵ.�E��fja��� ���F�W�U�H����䶟@=�L�o1=���=�S��w���$����=%= ����Ф��O�� �A��6�l�@�l�'�=@[A'���E�̱@h��F��*?�K[ٞ�{�l�3?��+�c���V2?B�/�?Tɉ��ZZƭ�:��ɂ�z
}��E��7�[��ÅJ���bL�0���u8(+C���O�v��2�Ǵ޷V�"�TH���1}s$�]�ǽ�gD��X���p?������nh���6���0R�9�=�h?&���J����C����G�K�B%�C($��Q�0U��w�+��]Mݷ:�V����5��D����GT�p�*���ӗp{�$ܣ�����-������Q�1Sx;��@��5��p7ci���D���aR�̬#"d�.3LZg������S��`��Y�K�ʧ4�0��-g}��֥Mh�c��\�m��o"(9�S���6|��;�0tT�s�l�AA��뉀K�\��v�O���� ���,����!�ٌ��/a׻{�A�3�[�#����%��q����<��Qo���t�߽K�>~�������.�'nHۤgF�:2~�G������ÎC#$���p�Vj��	Ȗ�S��I��Y�=�ꓨ����s��`^M�g�p�=S�֨.�ח�����P��'-�T�DGѭ�(j�o���a��A��+6ٓLr���m��O�S��ْZ��'��+9	��:��yǇq��M#`���Џtt��8��ɘ�Mg`�,�=v�ݮ/G��]��<�0le[|\�����J��^'bT���N�1�`�Z��|���g(���5F`sŷ�o[�cS7C��9��|J�2A*�e��H����S�ёz���ϱ���S�B��h],����h�a�����͑�!�M�U4+�����j�~ZE����S��ŉ��x�貲 $�|�7#��O��P����D�D�2P& ��I��`-��~�[���ꭈµ�K����I��Yvl"p��j�1���n|�?�u;�؋,�&�-�;⥮^x���H�hWuO�1$Ц��o6w�-�9�m`�(�V��h�1��?�Q=#�cQ�ul���5\�K��I���)�֦�a�)�	��-dc�qF�hތ؊���?]��z�<�L�ȴ�]j9M����p��U�N}>=|Դϩ��ApT�Bm@�!x9 ���e0�W�6��(Ԑ�G͂�(���˱AJ$vgMk����Ŗ�	�gI ��-��1��|i~ �IV�S��*��2������r�O;����i/[y��/T�x�ٔ�JV�@���~�'���?���{�e;;bS5e�t�o�%{�8���]��h�<��ȇ�v�_Ĭ��ZM�����,��^���%aW����/�d(s�&¨�7���j�jsa�FU�d�5>��:2�Vr�l[��%�a�����E��GJ�~/��z�@L\\�E�m��G=	uIy����|��x��OH�X�$'u�r��s J��kxX�z���t�3[4Tp��|0��} 8��Y�S.���S��]���j���gg��/����x��"���qd�%�������9�%��u����(kd�1r��Jz�Co�@)H��3�N"�8����Y��0�@Ǖ����7y_���xǬH�����E@5�����ە� Rf���F}�퇫�������
��'�|�K���!)��� ���$�vx�y� Q��M�����x�Y��ƪ})���1��܌>c����~�κ����Æ�<ɟȖ�]�����{0��p�S���@��ŠG�N��W7 ����̒�y��{b"���R`�c��G�#�_����������C*�ʷ��ufT���1�C����	�Kd+d�s�G[q��ѝ�3[��w�����@0����m��&�=@������V!�AY�'�e˵�6������
n���t��yI��V+�.v�#ǌ���҆e���N���4F ���6�C�v��MY�'��ϱBW�<����\�ILu�.}�'>��xi���ÍX-�t�hN>.��t�4���j}��y������㬸�=+�h�.Y��T]Cz��'�����փ�e��O⎐CG�[���i�ҽ%���)�mxJ�|�Ee-��'�7��l���c���L<���"q�CW�����C{��>�'�%B�.�1��PY����Ky+�{���B����k�R&����M����ܕ3|?">X��t[|����Z�����ۺ	~�ӕ��noc�!�͝�������	AH��l�P���6�z����5<��bA��t��k��mk
��F^�.Fؐ-�b��a�n�O>�,��	�b���j$�x9��\��7
l�ö���I��2&�$��Sr�i�5z^�Y�����<��>I�:Q�|��׶�"��3�|��i�[E[����m���gl;��!U�(yܶu>��َ7⟫���}U[|�?�tc����rkP����	E9�-Z�ZȌ�R0 H�t��r�g���d�������)�'��Ep���&k
bP�������S�^��K4)��$��8iH%e{	E�!���1��ڢ�n�R��XOd��o��)|Pk�Vj>@1'�b),R���a�pH���3i|��Y�V��<�s؅sEჩE6ށ��i�-�Q�h��vUXg}�U���)�3��|��ٝ?R�d>ݍC�� %�u}]�9Le}��;9ܤ_�v�%��L��>7�д���@�<� Ӕ�ԃ�̰!ך�<�+�I�Wh|�����3=-lf�⌒bApm��(���0�