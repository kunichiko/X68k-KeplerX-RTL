��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��5�������B���8���"���FE�Ҧ�@�Q\_������C]���5��1)2���� hڻ%pj�j��m���4 �w����4��O��� �P�˛����+���r\�8��s�;ۘ}�y���誛�I�e����-a�j��,C*��������~���>��75p�KcL�]�r��oՌ�I��r뎌 (��,H�grJ0�l���C-v��)���d�GFZ�bjU�zȱ%T��tz^'�kC0��&<ֺ�X��2I`})}�#���(`�p6V�I�䳥�a���#�]n�ù�ɚ�y pcY�0B� 0�Z��=�?�������V� k|%O�ܰ8��7i}kv���r(�F��%)�#Ua�����5�l�ZY��#�0`��:�u0�ĩ�ʩo:j�"�j<���i�s�P7W�0N;�~'iT�F��:�h'ne�r]i�`�����0�HK~�V�F>�P�@��n�wgTޔ`Ɔ�����R��`Dz�!*��3B�6�"ֹ�j���%r\�s�b��( ?�PH��{�1��{4%z]��O`�����X*��R��?O1M�=[F8�"e�*W��K;a-zt�"�� �f_u�^ �x��߀'��|�`���)�@h�j�Z�=N�1����!��Ѵ2���>5���:"�$�s!RhD���Pg����`ˑ�פc�$B/+d��)9��9󐢐ͬ�=4�Զ��u�k'�]��d�ԖDl��~O�{�5������P�`y�%�jx�:#���[��V�y��(���}؏�&ӓ�6v�k|��P��Ǭ ����Q�>,��bb���
����ms <�Y�5)��6�|n�JLO+�f�+�	'�*q�-�:
�揟���Fg0�������]�N%I�aZi��ԟq@&��O���RE؉X�NT�Ⱥv�K������q������@�d�U
!D(7U;e�I� �R[���x#j������y���ߚ�R��?�@�!A[b�{�����G�iBU�䐅������`�0��v}B���/UU^�>�O͖;~*��P՝ZT���n���&j~b@�VB:�7���!����`5'���OG/cfk�~��������)�Mw�u�2eQ�����s�_�e��I������E[�L�A9���pUt���|e��b��/���?��,8ᛳ<�D�D��<�GegT����9�&Oc~�47�x�@���P��F����D�s�Rj,��R���*�*{qk�S������#��%u�g�=��iT7����V���޲9��I�U&w#�ꅨ���̽�� ��o"��]��~�� Xy�%�kĥ	��uy�Ft���h�J��!��5�66����Y!�J�1=m��x���V��!����j��E]�L��.) �K�/�G��xQ���>�_篖��W��+9'$�Ŏz2��v���=�G���;G$�:�m�>u��,�C4@�<eF�4u'H�Wa�e�m�t��v�����NKYH�H3C�_ar�6j���-���H��,�x��v���݃\�	J���X�t\�6�]���0 �t
���X�w�ܤ�D����8����6�X,[�l"Mcn�z{]�{*���&���F�=�$j\G=���rZ�)����dD+@27�#���a(t���rԛ��\�)�;~��6<���$D�P����s%��j< <įW�\�[�}�c+�*�㪀:�d:6}޲݄�j��*?N�{.�0Y��H���I���2qx�P�B��� ���C�Ⱦ���D8`p�5��fu�WT �|��F�ōDx�g�31����¢�S�w?���B'�` ��T���a#��������kne�Fޕ=�R~s���8��p��54���CS�\�--���]>�ӛ���P�Fzmūg�@:n��nL":�2���:wH@�@H�Q�4�u�h�:���c���-���\쯔�$r��S�mx"��6וǞ.MF�[A_d�q����t��(�����(��	�>��&�v�Ǵ�;�r������G����ȕ(j���-a�B$�z��mo�.}3 �A�h�Zw�"��D2���c���n�%���h�m����뉀��G��I`���Ȏ񀓧��n u�	��g�陁�xU�ӱ�Eɂg��j�JG��r�EN �f�Z��R����K-ϥ��f{��O�]﷣�&��������_5�;����4An�MqH���-�F����ՙ��+,���?��:;�}�x�cT��'�A��C5��fzO��{��c9y��c�m(�*�G����}v���`[��3E �����0�5ַ�=+�_:cE�AG}���|�T��9��ߗh��#�G~�:�m��o�"�9�)�G�Q.�����/��+��'�'���o�K���k��lPw#�[hzv������qG�|8ˣ�a5��e�����|:���&6��O6T���g�)H?�p�T�g�&n�\�i,y{�:�k9��;�y� NdsBV�*�P�=M�W�h.�gc�44�8��V�������Y��;����)h'�1ʲ��<�i�L��`�F�����үK�G�nD�O�򺌒Ovs���uU?8¡��kHܯZ$��DI�j�
7%���cT}�n�C��/YR~�k�'��D>,W~X���Q�bX��j��/l��[���QM�sSC�D�:�j�9^��j�Sٌ*]c����S"O�����*9��c�UH�S>�q�c�ۮ�6�M'�!�L���!�nmٳ���Ժ���~�\�D�~Lڲ�뮛� v��TL�p�!WCG��N#
�]U����x�fz�7���$A�j�B���|�s�l��~zq7�cX��)r~#�@Q�2�N�e�:�hƽvk8��)��Vq���՚]�ʕ�����&!\�?��K�K0�d�������Y�o��O���E9�qQL����ն��4�����c�$�9=?I�u-�i&ԟ��{��e�ʳ�;?���a�:��&S|;C���HQ\C_�v���'>U=cA Zg�U�q9p��4��6L�?�{�H����F���K����M ��������&o�2������K~0��ZM��2�!>��o���e+�\���P�L�,�`v������DO|P4g��� ��]"��`1<S�-�%躳OB��
]��k�FNG�� x�RG�5u�-,��(���� �I}���ө���p��Pwl��Z5�E�5[`����ts���^�9���rՋ�����fJ��4���.���;S%8�Y�g�M�a�6��F�Z���!��L�۵�	g��1�ߘ3�͎���"+z��$�g�A^���`�w@nN�yD|� "���
�y�3�`@?7P�������z�=C01V����Q�1�N7D;�Ԣ��q���d�/�Ώ�����W䯘m���g�45��i���-)L F�F�7 z��(Y"�� �a��ޖ��z�\�������d��jAg����[m�I�!Wr���HxyN0DA46��[�~2�q�	>W��z�#Fp�`�p�����>��h�=7W�`+��`z�޽���P����sjd���ŻC��ot�^d�S7 �:�+O&,�O�z�/�h#�շ����_�RZ��^~�g,�{�E���2�F���r�;�DqyLc��M���+P���Ja[�a戼L��~D�[�j�,�N�j岔�6��c0%���g�j��^mB��������v��8��5�9{�rRk"�#�K��8��`�������=ܗq��D�r3<���?Y��k�=`�Yj�0�y�+������W�X��TmO��%�b���hQ&6o�"�c��z���+U���xME�=��uc�
�Zx�P��ʂ��n_���>�'����n�z4��k*�b����#�jͣw�n#�˩�r���pP#�8"oO-Q5ķ@�9���bؿ�	�O|�(��K	=�-'���D^4-Ce{�J�6���� w��d!�R��C��Nw)!�����p�m ٣ox�O����Z�2bV� ���iQ��3� ���:�M�mL�L�}绾R�{.��(~p���I�lp.D�JŊyј�h1��#�(p�`�q�	��Ժ�9� ���%Z?v�Y���Γ���!bL��YR���7��sOT)��*���9�$1�U����.�J�mq]t�[�~*!d�z�qys޼�
~K3Z2�>wdd�c�`�h�?��zɅ��g�qG<�+�-��L'_s��Q�* ��v�-�~��!�X(��R�{��ttmM��e�Ee��V�e���+�Jni�P��UK6Z�s�İ0��F~��<4�Z�����7]�V�%2@X��e����V���t�B�iR�Я���	���$̀��q�����2����7�h01�q����D�j��%W*���Xlup'�( �*�:��郮�ʘ%ˆ����/�������%�=�k�b͌Q�'� ?[G��\�0f�c�_��\�v������_�4�,�|���:�(5ǟ�#�Pc��SdP�n������S,L��Vm�C�?Ё
��q�{�m�1�(K��+����[�)��d�U'H��� ���=�q��D��^g�%��kC�f�2�}vP�����UoԄ<e]�Q���\cEϮ&oύ =f�_ѝ��{��Z5^e����V6w#W����3���j��.��^����@�<�����C'i��Y�X��tL�}ֽ�W�Б��ÒAz�>���Z~*Q�B[U��l�WsG%���C�$ie/P��·��^h�u�
�|����9bN
VdKØך�r�;�e��̞��k彚j�m���ƜQ�O�ޣ<���_��dr��JM0�,ӯv�Ǘ�v�h �]�8�G��9�l4�H�ܵ�bn�l��;'�z*qy�p�+��1eH����������G�H|r�CZ1b�Ę:� ���tz�cN��_��{��z��͎�)xcg�ԟү(4(vrB�̊��E���8�X�U�ۀiǑ���+��.�����A>&�4m�6.�hti��B|Ug6�Mw4��,�����Ox���6[G$�\��=H�/Z��r��߂̅�n)=si�P(��0�*w��Xe�w��U��S��8hHa����z���ecε&`��y�b@S���6��������}?ܿ�:@�e2�V�yH>ݛ¯�L�n�gKn`Wt����=a�1���j��a��q&�>Z^H�yXE���Fơ�[�lS�Ǫ"�����$p��ؚD܂���l#�.7%�c�.|�g�B��ş?����M�,�;�ss��TN�ڸ�(C�q<t��q@�ML�ɧ�a�P���������(�E*�l-'ՙ�<�(7����SfB�~�U�a��pK��Fu~o��d�G���U��k�aj�����9�TR�&���f��2\�T	�$��ҲP�?�j�Z ?_ُ���z?��%�����:�i/1�3�V�j?�����'�ҩ��R}��%�!�_�+���V�����N�M!���$]�9����B�z�E�Y7�d�_.��Ӷ����s'ҨA�,+`�