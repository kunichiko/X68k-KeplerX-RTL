��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D����gP�������������44��Pg��w�k�n�L�t�=�ʠ̲J�=�	�$tG�讧��p,��sC��Xu�_ S�	��mZK�qnu�*u"ǋ<�L*�2S���!��i�އh���
������)�=k��l��hx��I��} ���l��CaoK^G����F�HE���}�-���8���C��)�6v��q+���BɃ״��0�Ўl���Ax�`93Di�j�]��0x��uHo8ȁ�h�+���]�,L��uS��|�>5��9�8>�U̒ �|�o=���{�
'�[	��ԄgI.��Rs���Z�GݲB�_/h�_g�ˢGmYAa/E���,Ӥ`�΁b�d�@��+
��kz<ˤ(�w����0C݊��L87�C��������z��H�w��ڻJ�:>A��>I�B	�KW�-H��
 �ѶJ��;�\�16Ji�,�z}�:d�9E��_����Z���o-�[Ɯ��F$v�KG�%Z�:�oA4w�)[����:��z�X�o=B�e|�_2��ͰUSo����I#ظu��#x	oC}�v�%����KBU�2 p3 e�+�0ʝ��l�;$랉�A��t�h�?\�<��d"]���xuB�@3�{��e40/���GC��������ھΛ�HWR4��M�q��q��x�Gf�5�AW@{�-��LX�d��փ��Z�$�|�t��u�z(t�]7C�ua�Q�t��>l̘�9qaD���5:Ee��LsQ�����yEE����c��!�	B���IM:쐩���V���@���0��h�J�CX������7EC6���E9�c��"�Cޑ�.9䪙�Z�f�!3Ds^��d6з>m	���n�Y+�v��-#r��\'�;��o��4�_N��I	Y��>�N`E�C���7���9FkJU��v����Ga� �5��_�g�ѝ�k�
�h��ÃI������7Xΰ,?eVj1A[�^���/�@�I���sV̟r�<�7�m)�[���Ĉ,yz��k"/��Lh1T���(����b�\7���i��C�������/�����x�c6;��Y��ҟ.#�PJ��.]G:tD����⮾�5��HT�^��z��KG��!¨��E���R;���$�9刿�ds0��+O�O�[3xW���U��He�Ǵ�|[X���u+�'g�`�]ņ e�}���i+�?uN�`�~�"��դ�y��f��b�:�L,L2R�Ŏ�˓�F����\�IY<05�t�����_O�6��K[!Jޜ>4nag��+Zv�-֢p7���K;������O# �Q��ɤ�@�i���G��CZ {��A8ѭ����Ȭ"��P�_	�^�����a�{J���^�(���St���g���#��JƏ�����d��y�j���]%V��3bCm�� ��bi�=�t�S���l��o�H0���u�*��j�ZɃ�Jy���l_��"��@�񊷵Ӂ:d�D^Ek�5Д��]�����K�6KxLA^��EYHu�<��-\��DAl�[�����TT��4�C7�{����M(iE��������5��:TR��CG4 ���w0�XXLx,������焙.k��}���ꋀ�y<@jL�'�_P�G��!�x����y=�`���꧀d�@�OI���%����O�b�j��N~�-�3�5��ZG���t�}i����+qcr�	�NY_UwVd��\�ST�Dއp<@V#Q��H��9�S�^��?a����׭ըr%>%����GnIe���e?ND�������Zm��c�u#4������Z�a�i8q�f���"�����<��C�/�B�h�cY�����g����F�������:���3� jK�SF����Y����.���os�Hud�|����E�
s����n�h!OϞ�Js��k��/��Us&�g���|���5�xټpQ��=j�fc��ʠQU��/���tkDê7������� �[8���V�����vC����%w0��k8ѡ�E�:� 	fw��+e�D��`S���ɣ@B ��;C6+�.h���
��{�y�e��r�K�/����7�aFiU��B���4�l��?�wr�j1\�p���c)��D�����H�φ�E*�������'YE�\���Ռ9�7y=^�qT���R-
&�ir���_�$2�u��ħ�1Nz�2&�m&��t<����r�5��a���(�ad��Ly'F�(�1.k]*�s��^:�1�ǚ_�)����3Ã�������~�=����t�U�%�w� �-�4��Ȧ��
�ʂ��&���a�<) r� Ӕ=��$�6����$�@���QÒ�����|qj�~��K��Eb�~��{]h���@)���-�c����
_����xFK�h���ͥe�]�1o�}S���I��� S�!��Ʌ��EE�{�V{qh\O}+���q�� PH�
3�������F��e��3�G9����|K.g	 9p0*�9	�G����ZȬ����֭>}�}������A� 5u��Z�\th�#�2<P1.d��uY�><S�#�F�S���$�G�6���5�%��Llw�j�.t��O/���6
�54@U9��.���v�q�S/|YI������;��E�U�U6����I,���d5��0A�/� �=��/3�|5?�R����u~h�(���2�z�»s�o:��/���Ӿ9O!��>'�d�BH�����m[��x�t�T^Ͽ��Ҡ%�F���]�R>�s^��$���oS�"�I��!�+|c�
|�
��(��)�X�i�b�n��L�@r`߼
��E�T����}�-�}M �X<Lr8��V�7S�ٱ@|O��D��`��`T��p������
M@�e�����6���S�	�b��1�o�����Pmfj��88�X��A���[�������P��r��XjX5�R��sA4Z�^�bʿ���_�aC���)���n�$ �KQ��f+M��݄��I^��[��l��g"�}ۀ7��r��4v/�3a�j��tW}88TP�"�m���I���j>�p�f��l褛�A��h�5�0�~L��,�d�,	ȷ�>M��x��Qo]Θ�؛��!g1X>Jʵ{x�q�9���N��u�@�b:0r�چ�\�+%�z<�ҚZh���0S�!C���������Af�2��GuY��Ob�7��	��pT2�NI"b��9*�eK��[�]�w��^�/L�\!5]'Wm�n�ˍHE�dL��4d����<B�[�-Z���I��caD���E�&�"���j�I^L�ʤ``!�/�U�8~�����Fl�:?�B�Ft��E}b���z �{���-@A��O�)�\$MG��°���ۏh�OL�Hb?~,ǖ<��A+{NeҌ'Pt���/�y��/
��f���C�N1-�,��x������ 2kBN����<?�e��i�v3�Q!���:�O>Ť�Tך��~�w�q`A�m��3��.N	ݞ����J���\b��M:�f�,|O�L�J�^�h�� M�bJ�u�1vN��#c3�X�����=�e2���}��8�/k�2=u|��{)Ԃ����YU�Ǌ�^�`�D�3�����m�Fi�s��U�Fs\������� ���-36�CG�=���`�$=�����M�V+�{�[e�`a�˿>��o��X��'yd�S�ڢ}�,�3�c��w��`-�J�;4�����ƿ�3��w���-�Z�..���G]��gÿy� ��hʐ'��,
�ΔFy�< ��;�p}�Ԁ>�="$��?�{�����	�ӟ����Ei{)�+?%�h6��E��| ���� �����Vc��L��Y-��:�
Ȣ�)	�*?���RB�� �
��d��\\ׁ���ʉ ���C�>9�a�k˲���C��tX�J�*YZ�p�\��Z�&���뇍s��R9�EZ�$�Mk"�P>�SM*�k��1T�Vm�0,��ܛ/�zj	�g����Ee�p͡�f�>,��_�L�ύ\�$O�H� �Ԥ��V7Q��%�SV������L>���]�t@B�E{�m`���P&tt/>b�s��sW�%��&D��*޵�.Bӽ����,�B�0���L�!��2�жr�0��!(�A��nf^�c�j�l@F6՛>��E��uܘ3��Uh*�O[KZ��d$+��R���=���o7,w��`����m� 0������c{�iFf-XJ��J�BTQ7XĞ�h?`�K����l�s5,����5�^�����7gI�K��vqX��ET� ����l���԰���XPW,��&<%�#g��z�Ӑ;�t �N� i�JC��~vN/�V���E�7gPނG�M�����2}�?7~T��N��4z��,��@�1���fC�����C(�O�DۜOS�	�<��*x.ޜ'�-�����Q����	U{�-z%dn&t�:�yl�:�ZF�/٠R����@�f@�k�����I	0�R%�_��
����ҟ� ��>6���q�J���������\��(,GF 5�ʕ]o�O��ֆ��#u���)��qs��2Ќeʂ�p�ґ9��_a��'1�K�'c�B��t��yֳIE�>v
S6�X'��\��{_�x��`Q�s	A�d��N�����ҏ��I3��3�)g"G�$lI>�z�_����l�� :�����\&�yc,��G��r�'�rk�����`�~�ţ�p����bV/Mkϫ�4KIÝ7/�]P���L��Y���g�O7.�I>*]�}�>����b��4���D.���wmG����^���+�a�s��A��7� ��u@R��J2�H#̍O�+��7&V����{3^1Vx=~�7COR�๎6�)��(���{*Kk~�:�
b���oj�f�[�ngd
�=�X~��?����@�������˝[#iѴC+���>��#>����s���q�Yr@�`�> �O��x��>�ęm#h���%�H�n
�y����I��@�Ns�?��a��tE��KR=�u=B���%
��Ć���2�B,b�2��/��]�bs>QD���v`�*���PN�j�L��Fl�2�5[{>�TB��;ʤ��{:y�4��a8V���5��y65��sfy	1G���Zy+F,�B�y���Xz�訸�1e&���v@��(I*���z�+�r+�Wl��t�|��ӷ�Rǀ_=�]Z^JP£�_۬_��/�u%��K�JӋW��u�t�*y'"S��5��¬��!���v��{��P����2�[� *[��|)[��r��b��{��� ���U�z�5��:G�K��b���)�z�]�Q�#�c[@8��I ��d�����3��\8��p[����ѵk��9{ZӋ��9�ן��`@�2�*�L6�ѭwz���<v�<}��!v=q�]����T��햭O�."7,^ŧ��F��[�*T[߆�3&��F��������a��taUzh�?�l�� +Ĥ��p|�w� pg�^���5����c�S��)R|8mt�V���z�_����w�� �)Q淴�l=��ݹN�ti��6L"����
���,���#;W6tΑ�Z�E8>�Ƥ�+��5t�t�W!f�m�AG�;�YR��O|�{���#��^5�X�+<����q��0�u�r1�(+�/��D�L�΅k#=a�����a��w��~���Z�Ս}8*0E�?�i<)޺­��m�	�#'�ƭI�yDT�$�<8�.�ra��{�5/�o������w1������w�a.,}��{��ۙ�������:Ქv0&�Fớ��Kx��EH��������P@Z����4>�u-?m	a�
��k�-ɳBJo�z�F�P����i^�ͧ�=H���jx:)/��l�:1��O�~�O�8�Z�B�sꪍ�B#�_uz��Z�6@��50y��ò�3l�)�Rj�4�'=a��� H��?�Ű�%���;[���8���|��D����ر���C����$��nq	6�\eb������C��s�=�N�n]������wh.��.Ėo�H ����EI��K�i뭹Y�� G=,Nz����7���%iM�G�W���#��eiP��T�9gr
�Ŋva�|�@���#眬]�0����I�{}��˛�����B��z��G�D�Pd����Y�[ if2$@���@�.�ן�����hc}���8鞑�-�P|=�)� S�(ʂ}W��0�EX��y&�')F��B�ܴ�%��q���kv�?\ZA�[8��+�`8V��68E�o�@~4�4�ʛϖ�7��L��˂���j(��:=�
l���|�B�����"�O�vYY�E���?F�Y�L�R��74}��<��wG���\��v'�J�q?umE��g�,�*L?;�?��v�ð�M�1���v·FwV��⯁�_B~���W��\�6%lE����5�ٵB�>��������J�>رB�7�<��;d�$��+X���>-PK����l�B�7�y�,�a������Q���$��g�4�ۏ��E�G�z��6��"�#M��1{Y`�X��u�K�|�#w���̽�b���߄�]{�tf��wd�o*Ա�y���/�5�o:d��ƨ�L���)k�iv����>������|
��&Z�^�I���G�:a���Ma=K!+������ew֌q�1ʬ?�~��j��i[�U����Ka
�4^��}t������Ж��g�� �+�w�5̏fB��"Cs���k^l���<yM|{�E�%�y@	��/�����S��[.a)�&�p��t���;�����o�0m	��M:N7Lm����p�C����lVN<����Q�/X�����{�<j�O��ރuad�e%y�eS ��t>���
.��Y���5��jKd$���j�
g� }̦�KJ�0B���/3�NZw�'޹;�����0���]�/T�l�zq�6h_��[��dnc��b���IKm�ͱi� _z�g,[Pә�P��Hw�����0��P�f��k7�<��֯#��5���8��D޶�޿��Ԡ(�L�hH��=�IkG��()xe��K�G;~+�9c�S�K��&��_u^���p���{I�����-7�ON`�
=h����A��N���dO4�P�+O#aw�j�@*��{��7�o1��Y�l���r�ڠ\�!���P�̼�����z�#�3�'�h�iG�X�ퟝ�-�vw�3>Vc�g��r!���?V��N��@0�F����O6N��|�������9�Gy����e�*j�dH��_
��`�?2ܜ]>>�el��n��C�Wmw�ddך%�[���?�@��sm�� V��咣����e\���d���e�be��>-< R�Ȯ-���E)�P�K �/)u!MZQi���:�e��B�]��+t*b�p���I��T��R��*ZD���7&6l?�E�!����;�`�����9�?�����*���"eU%����8�!3�����ъyx$��'�N���̓CG�<%�;�Iմ��u�B.��e��B��x�����e�� ����'-(�����/pe�.�5��Na����Bo�i��P�Y"@�O�
�2I��B6�������wD��&�z�K����6�)Mg�S�7��Q��Q��m c�TY�� a"iJ�kds���68%_��fe��M�����q�쁣/-����\��r7I�����WB��w���V6�?�Yद�j0%�W�.ډt=�ؓ����)E5��f��c���,R=�Pp�B�jL�1�,��V�=�r���8Y��@�3��x��/�[��o�R�6��賚O��z�?����w*��UJx[N`d���C�GWP��y�S�8�.�I���1;�^�f��@�I��W��ڔ����#m�m	:�S%J�0���N�N�����9�.�YU��?���Y#&vE��ly��=iZ[.q'�D��4����������>�X��&��G_�X��͗Oy���{�(�x�����'b& �/�Dty{F�GVH@�BPP^�hx���s���'���.Nh��� r]��D�C�?=�ZB�\�Ƥ��T1�u#�{�E~"e_����3$!��p�c���D:<�|;% ��V:��$�P3�?����M���������Z��9��P�>/2��kK�ˉ�U��ґ95 ߳�ݽd��`yO�S�� �O������ɑ����n�0	�c6����5xN1�e��"�`��p��Q�e��ۀ|�f�B<�V��|ҙ��Q:����RF�3>�C��/��s�dA�VxhL���s7�4�[�~9ؘ�X/���R_�"C����ڟ�+½�HԚ�J��v����j6X��/��$u��\U�iC~�y�L1TL���9�����2�4%�Ύ/�U1��D�О��lod�q&�x����&m܎��fE6!�1<�[@\)�U%r���+F���ϟʺ�M>$C"�ن�#R�&5~�#��P�fw­~.t��I��3�M�&)���Y$�e���F���Nz�:!�tF�-f��G.�w����!�1��֜�8���A�0��QO:�z2~��_�U8=����{Z�u�{�:�F�Y!(�"�7���|np1�߀\�򥢆��qQ�k���*�2�[�Ձ��2��T���*�Ie^��* !|�[+z���w�JYC`�J�>�"*� ��2|��F�jЎ*9�BAwa�g����=��0��F�s���\ҫ栄�(�vb��	����Ӈeޛ�S=������'ܫ��G-�5�aW�v<7�0�:]��V��u����؃��s���L���#��(M����^�Ձ�j��פ��?�"챶�TtA��u3��[� ]�{�۠���T5�ƭ
��Jdhk�ר�^4��Z����U��n.��$9�\�VI'٤-J������X̛LDY����ু<m�W��IN��^B�`qZ��GB�g�iw�xܚ� ���~:c��Gl�^�*��uO}cZe���_��o��Y��y$LhKwSۢ��H��X�y�LD���E���LEoL�?@ 7l�_�����sÆf����,�[�9�r>���;ߋ���5�[��
g�]|�i�cV���.�MdL�O�]0���uNڦ��q�=���2�d</9�x!h��60�9�����r�������|?�A�AƘ��C>�;�EW���q,��"���i_I1�)./���e��K�����g��$��j�ՠh��������]��P��Y�V����#wE�s�Nx~�ٸ@C��'v�S�Ck�|62n������Z��v�	�k�:�]T�F��-�E���3�9���z�M`�]<�c�P�4�:@+b�q�i��!�&�1U�\3����8�)�����N��N�>�dQlm
H�N�����ic���,��$�܀�$}(�� ar��A1_�:�&�����6�zM�{Խ!��a7P���n�g8�S���>�n�5�5!WǓO̴\k�-�o�xt��z�t�����'�����z*$�s��4+�0�K�d.K+`�J�No�T6*w�k�܇�0��� �����dQu�UڮF��(UlrD�C���)�S-}�nw;�q����C�J�ؔq5)��rs��u�#y�%�п���~&����-�\�����b�^!���+�{�U�K}�QC]�`�ӗ�%x]�F�!	�w\V"��8�� E�4"��t�"R(��R6����Ö����Ȥ�E�Ts�`�H50�W � fSu> �Dl*�Va�c��f�u
|~��9��Æ��4��$�Y��Z��~,�m飍hdHS�n�"~C��t�� ���Ǔ�*��E��C��#���[K&o����q�=�f����y����vkV��i��D�Z8��h�r�Sh���	oO�y8*̥������o:w�mթ�o�p���|p9�UB��y͡V���0}�_U�S��~����-=��:2�E�/��I�#,�tP��^�G����T�L�G~��;)��e���1UѓU�d���Z��é�8�>ۡ��5J�Z=R,H7\*q���`5��D!Ȃ����I�X�����Vr���F�b:�[>g�B��M�$���\�RtX�4NFK�C�ձ�DT��C(Z��B/�JD�dlj���'�n�&��&����N�c4�^s�T�	�}Ĉm]+�:qFo
vF㖺B�"�mR�l�[������[^km�'��QQ䵥H�Z��2f�9�jQbB�6�K������It�Ҷ�L�H�}��_�aK2x�Xm�0��K�i� /ʥ�6�:��K���X��V�R�Y��8�3V�arO�9Ӕ����E�!+�F0cp���*��?�)�`�>+dPu�W��x.�"<�a�6��JOIe%V�i��.�͹Vd��7 ��Dd���c3�Q��u.j�7���Ni[�}K��8<	�B�+ͅ�l�w�L:X���!#%������׊���j�����;�����Ҥ���R�]pR�6���Y>�n���]���̐���f'}zy�h��ڬ��T��_/7��2n��.|��Se�r��TD2�����=�͉}�'�zQ��I�I]ƌ3��]b�Q)���X[*������8�ov=�Iu�������R�~��f�]JM�*w��#/̭�d+'N��u�$_�QX����.�� �[4T����u�s�D\�W$BR��ִ<.rn��p�2���)�a|�zܺf�kJ1P|T)3Vn��G���%�g���>EB�L]!�^�Il�*`�9"�n�<��4A�[��Ng��1�W,�в0���,��
q���P$5n���Ǌ}]eh0թ]�S �]�����h2��֜ܛF�lf:j���m�V��1�،#��+�a��7��	}�R��.��jB���u09���L�����!��9�d�xR4�_&չU��ʵ��uw=�m�M�����F��j��,�m(��bM8��.�.�-ʠ�%^�m�c�ںw��<ԡP�9��z�j#� MsI��Q��(x�Ċ���~G���Ms�tm��3oy��7�dj�����wr���i�(2|:�P�$�tt��*�7���d"��eMf��_B��ː�s�+��[_rHD'%��~e���gC&�]�b�����)㻫$��)����,�>�t3��d_#+u"R�&-�cC�^�#�53&��w���6Y�Q 9k7����!OP��T��؎Ep�^��گf�ZĈ��;4\�?���)ٯs��6�V���@��D݂�r-=�������A2�������D6(2�����Z� <�/܅��WB^*@@�$���77�%������ |-���֢$Z���k<��k�4���[��͇��L��]�%\hq+v�l�$�{��W�"o��'��|d�N�?�G��px�A,��,����<QG��t z���T
���p��<�c-^ S<I�$f� }��~+��rR)�q���wޣY8�;MYW�vn��<E���S5��e
�z��tl���v����&��n�QQ*K �f��2nNUbq>?q�g-���g�	���N�"
O ��t����+d_'�r��Z�(�x�u.��/���1E"�F���K�9��"'�:��#��Q!�:�i��AS>ρ���A���Y��B:�����m�N�L�/s�j|՘��}V�aR�n#�璨M�wC���(�4��������bH��jm�l�%(��,�8��]��Jͼɠ�@=�(n��+������ש��x�c�C ��h�3z,�(\��B=�r�����wz�aq��2���W�N���W|����8����=3��os�	���[��A_�\jvz�����jaX������R���2��+���b:e�bz��3�uN��b ]j���N�7D}T/m���Kqƴf�$^��p�XO��@�t�LQP{���t���ѻf�OQ"�&=KMO/m�;��&Zj����fj���p�B��Ên��|-`��k	:k��X�eq��7�H֏���G@k�o-�yǢ��+n��W�z�,K��]2ſ�z��yRId�މqy����Y���"��/' �Ŝ'x?Ϻ]��b�n�s��p�%�-�\�h>�n'��[Qލ 3�}�:��)�>��\�{
�gAuyO�a5 S��������旱�gJj�;�az	�"��ޠN<���$�F��&=&k�iXɜ��'{r��ϋw�=����3w6��4Q��O�ooU�����Ӌ�Efʶ&dƸ��w`��?��A۴�����Y;!u֥s���߯�Yv,�.P7ty�RtΆ�S)�k�J��;Fϊ��Q���xz�f���0S&2�YD���b�+Ԓ��z�ި���W��M�@�xg(pW����u��S���\��n��@BI����� ̎�����[�Y/�d�L�������Й"O��?G��y��6�4S�|F��n���2�%�4e�;��� )��g�jr���R�4�+���b����z���f�<�Ά!U�tE-�#�A�=BP�IN*��H~�����pOmC�]�#Ɠ��b	���K�sE"|�E�8�,_&�s��/��T�p��y�?�/��j���(��T�K�tB�v�<��+D�eG�������<�0�C�[H��ȡ�����I��{M��N�c\����Hq�՘+�ٰ|��Ỳ���$vnnU?!���L��tm����x�W���IUN�/:���� �$%�"���P9i�Ї�����;��Z���$���գ0��!�� S���aiTBܖyݬ2��
�I��ｿ�C��1oV���iWd�*s���!Ȇ۪�C'�� ��}c-Is���iL���#��s��3w�w�c0�XYC5Z�̊�qk�SW ����D���c&:X�:�"��1���n����2�B��eJ,eS��c8�lB�{�}�z�z�[!Y�D�*@yT��|�w�lɝ�0�_u�\�
���"�i�t����;]��<�x�B�4�mݨ�/�>�a�r9�^AL���w�p�
���>�TSjqx�HX��Q�Q�"���_&�B|�K� `��$�$W�hR��q�6s6O�������'���� ԣ� �x